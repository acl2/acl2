// SV - Symbolic Vector Hardware Analysis Framework
// Copyright (C) 2014-2015 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Sol Swords <sswords@centtech.com>



module spec (input logic [127:0] in,
	     output wire [127:0] out);

   parameter a = 10;
   parameter b = 12;
   parameter c = 16;
  logic [3:0] foo;
   assign foo[0] = in[1:0] == 0;
   assign foo[1] = in[1:0] == 1;
   assign foo[2] = in[1:0] == 2;
   assign foo[3] = in[1:0] == 3;

   parameter width=3;

  logic [3:0] bar;
   assign out = foo[0] ? $unsigned( (width+1)'(a)) :
		foo[1] ? $unsigned( (width+1)'(b)) :
		foo[2] ? $unsigned( (width+1)'(45)) :
		foo[3] ? $unsigned( (width+1)'(33)) :
		         $unsigned( (width+1)'(c));

   // assign out = bar;

endmodule
                 

   
