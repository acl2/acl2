module top (output topout, input topin);

  // Can't have a zero-ary not gate
  not();

endmodule
