module top ();

  // Can't have a zero-ary not gate
  not();

endmodule
