

module top (output topout, input topin);

  import pack::*; // package doesn't exist

endmodule
