// SVEX - Symbolic, Vector-Level Hardware Description Library
// Copyright (C) 2014 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Sol Swords <sswords@centtech.com>

module test ();

   localparam nCycles = 1024;

  reg [127:0] inputs [nCycles-1:0];
  reg [127:0] outputs [nCycles-1:0];

  reg [127:0] in;
  reg [127:0] out;

  reg clk;

   spec specinst (.*);


  integer i;
   initial begin
     $dumpfile("test.vcd");
     $dumpvars();
     clk = 0;
     $readmemb("inputs.data", inputs);
     for (i=0; i<nCycles; i++) begin
       in = inputs[i];
       #2;
       clk = 1;
       #5;
       clk = 0;
       #3;
       outputs[i] = out;
     end
     $writememb(`outfile, outputs);
   end
endmodule
