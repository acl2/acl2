module top ;

  genvar i;
  assign i = 0;  // oops, assignment to genvar?

endmodule
