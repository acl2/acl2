// SV - Symbolic Vector Hardware Analysis Framework
// Copyright (C) 2014-2015 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Sol Swords <sswords@centtech.com>

package S;
   localparam BB = 4;
endpackage // S

package P;
   parameter UB = 13;
endpackage

package U;
   import P::*;
  typedef logic [(S::BB)-1:0] b_t;
  typedef logic [UB-$bits(b_t)-2:0] u_t;
   localparam u_t aaa = 4'b0?00;
   localparam u_t bbb = 4'b0?01;
   localparam u_t ccc = 4'b1??1;
   localparam u_t ddd = 4'b1??0;
   localparam u_t eee = 4'b0?1?;
endpackage

package sd;
   localparam AB = 4;

   import U::u_t;

   function automatic [AB-1:0] g (u_t u);
     import U::*;
     unique casez (u)
       aaa : return 1;
       bbb : return 2;
       ccc : return 3;
       ddd : return 4;
       eee : return 5;
       default: return 'x;
     endcase // unique casez (u)
   endfunction // g
endpackage


module spec (input logic [127:0] in,
	     output logic [127:0] out);

   assign out = sd::g(in);

endmodule // spec

