// SV - Symbolic Vector Hardware Analysis Framework
// Copyright (C) 2014-2015 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Sol Swords <sswords@centtech.com>

module spec (input logic [127:0] in,
	     output logic [127:0] out);

  typedef struct {
    logic [3:0] a [1:0][3:0];
    logic [3:0] b [1:0][3:0];
  } mems;

   mems m;

  logic [1:0] indices [3:0];
  logic [3:0] vals [3:0];

   assign { vals[3], vals[2], vals[1], vals[0], indices[3], indices[2], indices[1], indices[0] } = in;


  int i [3:0];

   always_comb begin
     { m.a[0][3], m.a[0][2], m.a[0][1], m.a[0][0] } = '0;
     m.a[0][indices[0]] = vals[0];
   end

   always_comb begin
     { m.a[1][3], m.a[1][2], m.a[1][1], m.a[1][0] } = '0;
     m.a[1][indices[1]] = vals[1];
   end

   always_comb begin
     { m.b[0][3], m.b[0][2], m.b[0][1], m.b[0][0] } = '0;
     m.b[0][indices[2]] = vals[2];
   end

   always_comb begin
     { m.b[1][3], m.b[1][2], m.b[1][1], m.b[1][0] } = '0;
     m.b[1][indices[3]] = vals[3];
   end

   assign out = { m.b[1][3], m.b[1][2], m.b[1][1], m.b[1][0],
                  m.b[0][3], m.b[0][2], m.b[0][1], m.b[0][0],
                  m.a[1][3], m.a[1][2], m.a[1][1], m.a[1][0],
                  m.a[0][3], m.a[0][2], m.a[0][1], m.a[0][0] };


endmodule   
