module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
    endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
    endmodule


module DT_SB4_HC_64_64(
        input logic [63:0] IN1,
        input logic [63:0] IN2,
        output logic [127:0] result);
    
    
// Creating Partial Products 

    wire logic const1;
    assign const1 = 1'b1;
    
    // Signed Booth Radix-4 Partial Products Row 1
    wire logic select_e_0, select_ne_0, select_2x_0, tcomp0, select_n2x_0;
    assign select_e_0 = ((~ IN1[1]) & (IN1[0] ^ 1'b0));
    assign select_ne_0 = IN1[1] &  (IN1[0] ^ 1'b0);
    assign select_2x_0 = (~ IN1[1]) & IN1[0] & 1'b0;
    assign select_n2x_0 = IN1[1] & (~ IN1[0]) & (~ 1'b0);
    wire logic pp_0_0;
    assign pp_0_0 = (select_e_0 & IN2[0] | select_2x_0 & 1'b0 | select_n2x_0 & 1'b1 | select_ne_0 & (~ IN2[0])  );
    wire logic pp_0_1;
    assign pp_0_1 = (select_e_0 & IN2[1] | select_2x_0 & IN2[0] | select_n2x_0 & (~ IN2[0]) | select_ne_0 & (~ IN2[1])  );
    wire logic pp_0_2;
    assign pp_0_2 = (select_e_0 & IN2[2] | select_2x_0 & IN2[1] | select_n2x_0 & (~ IN2[1]) | select_ne_0 & (~ IN2[2])  );
    wire logic pp_0_3;
    assign pp_0_3 = (select_e_0 & IN2[3] | select_2x_0 & IN2[2] | select_n2x_0 & (~ IN2[2]) | select_ne_0 & (~ IN2[3])  );
    wire logic pp_0_4;
    assign pp_0_4 = (select_e_0 & IN2[4] | select_2x_0 & IN2[3] | select_n2x_0 & (~ IN2[3]) | select_ne_0 & (~ IN2[4])  );
    wire logic pp_0_5;
    assign pp_0_5 = (select_e_0 & IN2[5] | select_2x_0 & IN2[4] | select_n2x_0 & (~ IN2[4]) | select_ne_0 & (~ IN2[5])  );
    wire logic pp_0_6;
    assign pp_0_6 = (select_e_0 & IN2[6] | select_2x_0 & IN2[5] | select_n2x_0 & (~ IN2[5]) | select_ne_0 & (~ IN2[6])  );
    wire logic pp_0_7;
    assign pp_0_7 = (select_e_0 & IN2[7] | select_2x_0 & IN2[6] | select_n2x_0 & (~ IN2[6]) | select_ne_0 & (~ IN2[7])  );
    wire logic pp_0_8;
    assign pp_0_8 = (select_e_0 & IN2[8] | select_2x_0 & IN2[7] | select_n2x_0 & (~ IN2[7]) | select_ne_0 & (~ IN2[8])  );
    wire logic pp_0_9;
    assign pp_0_9 = (select_e_0 & IN2[9] | select_2x_0 & IN2[8] | select_n2x_0 & (~ IN2[8]) | select_ne_0 & (~ IN2[9])  );
    wire logic pp_0_10;
    assign pp_0_10 = (select_e_0 & IN2[10] | select_2x_0 & IN2[9] | select_n2x_0 & (~ IN2[9]) | select_ne_0 & (~ IN2[10])  );
    wire logic pp_0_11;
    assign pp_0_11 = (select_e_0 & IN2[11] | select_2x_0 & IN2[10] | select_n2x_0 & (~ IN2[10]) | select_ne_0 & (~ IN2[11])  );
    wire logic pp_0_12;
    assign pp_0_12 = (select_e_0 & IN2[12] | select_2x_0 & IN2[11] | select_n2x_0 & (~ IN2[11]) | select_ne_0 & (~ IN2[12])  );
    wire logic pp_0_13;
    assign pp_0_13 = (select_e_0 & IN2[13] | select_2x_0 & IN2[12] | select_n2x_0 & (~ IN2[12]) | select_ne_0 & (~ IN2[13])  );
    wire logic pp_0_14;
    assign pp_0_14 = (select_e_0 & IN2[14] | select_2x_0 & IN2[13] | select_n2x_0 & (~ IN2[13]) | select_ne_0 & (~ IN2[14])  );
    wire logic pp_0_15;
    assign pp_0_15 = (select_e_0 & IN2[15] | select_2x_0 & IN2[14] | select_n2x_0 & (~ IN2[14]) | select_ne_0 & (~ IN2[15])  );
    wire logic pp_0_16;
    assign pp_0_16 = (select_e_0 & IN2[16] | select_2x_0 & IN2[15] | select_n2x_0 & (~ IN2[15]) | select_ne_0 & (~ IN2[16])  );
    wire logic pp_0_17;
    assign pp_0_17 = (select_e_0 & IN2[17] | select_2x_0 & IN2[16] | select_n2x_0 & (~ IN2[16]) | select_ne_0 & (~ IN2[17])  );
    wire logic pp_0_18;
    assign pp_0_18 = (select_e_0 & IN2[18] | select_2x_0 & IN2[17] | select_n2x_0 & (~ IN2[17]) | select_ne_0 & (~ IN2[18])  );
    wire logic pp_0_19;
    assign pp_0_19 = (select_e_0 & IN2[19] | select_2x_0 & IN2[18] | select_n2x_0 & (~ IN2[18]) | select_ne_0 & (~ IN2[19])  );
    wire logic pp_0_20;
    assign pp_0_20 = (select_e_0 & IN2[20] | select_2x_0 & IN2[19] | select_n2x_0 & (~ IN2[19]) | select_ne_0 & (~ IN2[20])  );
    wire logic pp_0_21;
    assign pp_0_21 = (select_e_0 & IN2[21] | select_2x_0 & IN2[20] | select_n2x_0 & (~ IN2[20]) | select_ne_0 & (~ IN2[21])  );
    wire logic pp_0_22;
    assign pp_0_22 = (select_e_0 & IN2[22] | select_2x_0 & IN2[21] | select_n2x_0 & (~ IN2[21]) | select_ne_0 & (~ IN2[22])  );
    wire logic pp_0_23;
    assign pp_0_23 = (select_e_0 & IN2[23] | select_2x_0 & IN2[22] | select_n2x_0 & (~ IN2[22]) | select_ne_0 & (~ IN2[23])  );
    wire logic pp_0_24;
    assign pp_0_24 = (select_e_0 & IN2[24] | select_2x_0 & IN2[23] | select_n2x_0 & (~ IN2[23]) | select_ne_0 & (~ IN2[24])  );
    wire logic pp_0_25;
    assign pp_0_25 = (select_e_0 & IN2[25] | select_2x_0 & IN2[24] | select_n2x_0 & (~ IN2[24]) | select_ne_0 & (~ IN2[25])  );
    wire logic pp_0_26;
    assign pp_0_26 = (select_e_0 & IN2[26] | select_2x_0 & IN2[25] | select_n2x_0 & (~ IN2[25]) | select_ne_0 & (~ IN2[26])  );
    wire logic pp_0_27;
    assign pp_0_27 = (select_e_0 & IN2[27] | select_2x_0 & IN2[26] | select_n2x_0 & (~ IN2[26]) | select_ne_0 & (~ IN2[27])  );
    wire logic pp_0_28;
    assign pp_0_28 = (select_e_0 & IN2[28] | select_2x_0 & IN2[27] | select_n2x_0 & (~ IN2[27]) | select_ne_0 & (~ IN2[28])  );
    wire logic pp_0_29;
    assign pp_0_29 = (select_e_0 & IN2[29] | select_2x_0 & IN2[28] | select_n2x_0 & (~ IN2[28]) | select_ne_0 & (~ IN2[29])  );
    wire logic pp_0_30;
    assign pp_0_30 = (select_e_0 & IN2[30] | select_2x_0 & IN2[29] | select_n2x_0 & (~ IN2[29]) | select_ne_0 & (~ IN2[30])  );
    wire logic pp_0_31;
    assign pp_0_31 = (select_e_0 & IN2[31] | select_2x_0 & IN2[30] | select_n2x_0 & (~ IN2[30]) | select_ne_0 & (~ IN2[31])  );
    wire logic pp_0_32;
    assign pp_0_32 = (select_e_0 & IN2[32] | select_2x_0 & IN2[31] | select_n2x_0 & (~ IN2[31]) | select_ne_0 & (~ IN2[32])  );
    wire logic pp_0_33;
    assign pp_0_33 = (select_e_0 & IN2[33] | select_2x_0 & IN2[32] | select_n2x_0 & (~ IN2[32]) | select_ne_0 & (~ IN2[33])  );
    wire logic pp_0_34;
    assign pp_0_34 = (select_e_0 & IN2[34] | select_2x_0 & IN2[33] | select_n2x_0 & (~ IN2[33]) | select_ne_0 & (~ IN2[34])  );
    wire logic pp_0_35;
    assign pp_0_35 = (select_e_0 & IN2[35] | select_2x_0 & IN2[34] | select_n2x_0 & (~ IN2[34]) | select_ne_0 & (~ IN2[35])  );
    wire logic pp_0_36;
    assign pp_0_36 = (select_e_0 & IN2[36] | select_2x_0 & IN2[35] | select_n2x_0 & (~ IN2[35]) | select_ne_0 & (~ IN2[36])  );
    wire logic pp_0_37;
    assign pp_0_37 = (select_e_0 & IN2[37] | select_2x_0 & IN2[36] | select_n2x_0 & (~ IN2[36]) | select_ne_0 & (~ IN2[37])  );
    wire logic pp_0_38;
    assign pp_0_38 = (select_e_0 & IN2[38] | select_2x_0 & IN2[37] | select_n2x_0 & (~ IN2[37]) | select_ne_0 & (~ IN2[38])  );
    wire logic pp_0_39;
    assign pp_0_39 = (select_e_0 & IN2[39] | select_2x_0 & IN2[38] | select_n2x_0 & (~ IN2[38]) | select_ne_0 & (~ IN2[39])  );
    wire logic pp_0_40;
    assign pp_0_40 = (select_e_0 & IN2[40] | select_2x_0 & IN2[39] | select_n2x_0 & (~ IN2[39]) | select_ne_0 & (~ IN2[40])  );
    wire logic pp_0_41;
    assign pp_0_41 = (select_e_0 & IN2[41] | select_2x_0 & IN2[40] | select_n2x_0 & (~ IN2[40]) | select_ne_0 & (~ IN2[41])  );
    wire logic pp_0_42;
    assign pp_0_42 = (select_e_0 & IN2[42] | select_2x_0 & IN2[41] | select_n2x_0 & (~ IN2[41]) | select_ne_0 & (~ IN2[42])  );
    wire logic pp_0_43;
    assign pp_0_43 = (select_e_0 & IN2[43] | select_2x_0 & IN2[42] | select_n2x_0 & (~ IN2[42]) | select_ne_0 & (~ IN2[43])  );
    wire logic pp_0_44;
    assign pp_0_44 = (select_e_0 & IN2[44] | select_2x_0 & IN2[43] | select_n2x_0 & (~ IN2[43]) | select_ne_0 & (~ IN2[44])  );
    wire logic pp_0_45;
    assign pp_0_45 = (select_e_0 & IN2[45] | select_2x_0 & IN2[44] | select_n2x_0 & (~ IN2[44]) | select_ne_0 & (~ IN2[45])  );
    wire logic pp_0_46;
    assign pp_0_46 = (select_e_0 & IN2[46] | select_2x_0 & IN2[45] | select_n2x_0 & (~ IN2[45]) | select_ne_0 & (~ IN2[46])  );
    wire logic pp_0_47;
    assign pp_0_47 = (select_e_0 & IN2[47] | select_2x_0 & IN2[46] | select_n2x_0 & (~ IN2[46]) | select_ne_0 & (~ IN2[47])  );
    wire logic pp_0_48;
    assign pp_0_48 = (select_e_0 & IN2[48] | select_2x_0 & IN2[47] | select_n2x_0 & (~ IN2[47]) | select_ne_0 & (~ IN2[48])  );
    wire logic pp_0_49;
    assign pp_0_49 = (select_e_0 & IN2[49] | select_2x_0 & IN2[48] | select_n2x_0 & (~ IN2[48]) | select_ne_0 & (~ IN2[49])  );
    wire logic pp_0_50;
    assign pp_0_50 = (select_e_0 & IN2[50] | select_2x_0 & IN2[49] | select_n2x_0 & (~ IN2[49]) | select_ne_0 & (~ IN2[50])  );
    wire logic pp_0_51;
    assign pp_0_51 = (select_e_0 & IN2[51] | select_2x_0 & IN2[50] | select_n2x_0 & (~ IN2[50]) | select_ne_0 & (~ IN2[51])  );
    wire logic pp_0_52;
    assign pp_0_52 = (select_e_0 & IN2[52] | select_2x_0 & IN2[51] | select_n2x_0 & (~ IN2[51]) | select_ne_0 & (~ IN2[52])  );
    wire logic pp_0_53;
    assign pp_0_53 = (select_e_0 & IN2[53] | select_2x_0 & IN2[52] | select_n2x_0 & (~ IN2[52]) | select_ne_0 & (~ IN2[53])  );
    wire logic pp_0_54;
    assign pp_0_54 = (select_e_0 & IN2[54] | select_2x_0 & IN2[53] | select_n2x_0 & (~ IN2[53]) | select_ne_0 & (~ IN2[54])  );
    wire logic pp_0_55;
    assign pp_0_55 = (select_e_0 & IN2[55] | select_2x_0 & IN2[54] | select_n2x_0 & (~ IN2[54]) | select_ne_0 & (~ IN2[55])  );
    wire logic pp_0_56;
    assign pp_0_56 = (select_e_0 & IN2[56] | select_2x_0 & IN2[55] | select_n2x_0 & (~ IN2[55]) | select_ne_0 & (~ IN2[56])  );
    wire logic pp_0_57;
    assign pp_0_57 = (select_e_0 & IN2[57] | select_2x_0 & IN2[56] | select_n2x_0 & (~ IN2[56]) | select_ne_0 & (~ IN2[57])  );
    wire logic pp_0_58;
    assign pp_0_58 = (select_e_0 & IN2[58] | select_2x_0 & IN2[57] | select_n2x_0 & (~ IN2[57]) | select_ne_0 & (~ IN2[58])  );
    wire logic pp_0_59;
    assign pp_0_59 = (select_e_0 & IN2[59] | select_2x_0 & IN2[58] | select_n2x_0 & (~ IN2[58]) | select_ne_0 & (~ IN2[59])  );
    wire logic pp_0_60;
    assign pp_0_60 = (select_e_0 & IN2[60] | select_2x_0 & IN2[59] | select_n2x_0 & (~ IN2[59]) | select_ne_0 & (~ IN2[60])  );
    wire logic pp_0_61;
    assign pp_0_61 = (select_e_0 & IN2[61] | select_2x_0 & IN2[60] | select_n2x_0 & (~ IN2[60]) | select_ne_0 & (~ IN2[61])  );
    wire logic pp_0_62;
    assign pp_0_62 = (select_e_0 & IN2[62] | select_2x_0 & IN2[61] | select_n2x_0 & (~ IN2[61]) | select_ne_0 & (~ IN2[62])  );
    wire logic pp_0_63;
    assign pp_0_63 = (select_e_0 & IN2[63] | select_2x_0 & IN2[62] | select_n2x_0 & (~ IN2[62]) | select_ne_0 & (~ IN2[63])  );
    wire logic pp_0_64;
    assign pp_0_64 = (select_e_0 & IN2[63] | select_2x_0 & IN2[63] | select_n2x_0 & (~ IN2[63]) | select_ne_0 & (~ IN2[63])  );
    wire logic pp_0_65;
    assign pp_0_65 = ~ (select_e_0 & IN2[63] | select_2x_0 & IN2[63] | select_n2x_0 & (~ IN2[63]) | select_ne_0 & (~ IN2[63])  );
    assign tcomp0 = select_ne_0 | select_n2x_0;
    
    // Signed Booth Radix-4 Partial Products Row 2
    wire logic select_e_1, select_ne_1, select_2x_1, tcomp1, select_n2x_1;
    assign select_e_1 = ((~ IN1[3]) & (IN1[2] ^ IN1[1]));
    assign select_ne_1 = IN1[3] &  (IN1[2] ^ IN1[1]);
    assign select_2x_1 = (~ IN1[3]) & IN1[2] & IN1[1];
    assign select_n2x_1 = IN1[3] & (~ IN1[2]) & (~ IN1[1]);
    wire logic pp_1_0;
    assign pp_1_0 = (select_e_1 & IN2[0] | select_2x_1 & 1'b0 | select_n2x_1 & 1'b1 | select_ne_1 & (~ IN2[0])  );
    wire logic pp_1_1;
    assign pp_1_1 = (select_e_1 & IN2[1] | select_2x_1 & IN2[0] | select_n2x_1 & (~ IN2[0]) | select_ne_1 & (~ IN2[1])  );
    wire logic pp_1_2;
    assign pp_1_2 = (select_e_1 & IN2[2] | select_2x_1 & IN2[1] | select_n2x_1 & (~ IN2[1]) | select_ne_1 & (~ IN2[2])  );
    wire logic pp_1_3;
    assign pp_1_3 = (select_e_1 & IN2[3] | select_2x_1 & IN2[2] | select_n2x_1 & (~ IN2[2]) | select_ne_1 & (~ IN2[3])  );
    wire logic pp_1_4;
    assign pp_1_4 = (select_e_1 & IN2[4] | select_2x_1 & IN2[3] | select_n2x_1 & (~ IN2[3]) | select_ne_1 & (~ IN2[4])  );
    wire logic pp_1_5;
    assign pp_1_5 = (select_e_1 & IN2[5] | select_2x_1 & IN2[4] | select_n2x_1 & (~ IN2[4]) | select_ne_1 & (~ IN2[5])  );
    wire logic pp_1_6;
    assign pp_1_6 = (select_e_1 & IN2[6] | select_2x_1 & IN2[5] | select_n2x_1 & (~ IN2[5]) | select_ne_1 & (~ IN2[6])  );
    wire logic pp_1_7;
    assign pp_1_7 = (select_e_1 & IN2[7] | select_2x_1 & IN2[6] | select_n2x_1 & (~ IN2[6]) | select_ne_1 & (~ IN2[7])  );
    wire logic pp_1_8;
    assign pp_1_8 = (select_e_1 & IN2[8] | select_2x_1 & IN2[7] | select_n2x_1 & (~ IN2[7]) | select_ne_1 & (~ IN2[8])  );
    wire logic pp_1_9;
    assign pp_1_9 = (select_e_1 & IN2[9] | select_2x_1 & IN2[8] | select_n2x_1 & (~ IN2[8]) | select_ne_1 & (~ IN2[9])  );
    wire logic pp_1_10;
    assign pp_1_10 = (select_e_1 & IN2[10] | select_2x_1 & IN2[9] | select_n2x_1 & (~ IN2[9]) | select_ne_1 & (~ IN2[10])  );
    wire logic pp_1_11;
    assign pp_1_11 = (select_e_1 & IN2[11] | select_2x_1 & IN2[10] | select_n2x_1 & (~ IN2[10]) | select_ne_1 & (~ IN2[11])  );
    wire logic pp_1_12;
    assign pp_1_12 = (select_e_1 & IN2[12] | select_2x_1 & IN2[11] | select_n2x_1 & (~ IN2[11]) | select_ne_1 & (~ IN2[12])  );
    wire logic pp_1_13;
    assign pp_1_13 = (select_e_1 & IN2[13] | select_2x_1 & IN2[12] | select_n2x_1 & (~ IN2[12]) | select_ne_1 & (~ IN2[13])  );
    wire logic pp_1_14;
    assign pp_1_14 = (select_e_1 & IN2[14] | select_2x_1 & IN2[13] | select_n2x_1 & (~ IN2[13]) | select_ne_1 & (~ IN2[14])  );
    wire logic pp_1_15;
    assign pp_1_15 = (select_e_1 & IN2[15] | select_2x_1 & IN2[14] | select_n2x_1 & (~ IN2[14]) | select_ne_1 & (~ IN2[15])  );
    wire logic pp_1_16;
    assign pp_1_16 = (select_e_1 & IN2[16] | select_2x_1 & IN2[15] | select_n2x_1 & (~ IN2[15]) | select_ne_1 & (~ IN2[16])  );
    wire logic pp_1_17;
    assign pp_1_17 = (select_e_1 & IN2[17] | select_2x_1 & IN2[16] | select_n2x_1 & (~ IN2[16]) | select_ne_1 & (~ IN2[17])  );
    wire logic pp_1_18;
    assign pp_1_18 = (select_e_1 & IN2[18] | select_2x_1 & IN2[17] | select_n2x_1 & (~ IN2[17]) | select_ne_1 & (~ IN2[18])  );
    wire logic pp_1_19;
    assign pp_1_19 = (select_e_1 & IN2[19] | select_2x_1 & IN2[18] | select_n2x_1 & (~ IN2[18]) | select_ne_1 & (~ IN2[19])  );
    wire logic pp_1_20;
    assign pp_1_20 = (select_e_1 & IN2[20] | select_2x_1 & IN2[19] | select_n2x_1 & (~ IN2[19]) | select_ne_1 & (~ IN2[20])  );
    wire logic pp_1_21;
    assign pp_1_21 = (select_e_1 & IN2[21] | select_2x_1 & IN2[20] | select_n2x_1 & (~ IN2[20]) | select_ne_1 & (~ IN2[21])  );
    wire logic pp_1_22;
    assign pp_1_22 = (select_e_1 & IN2[22] | select_2x_1 & IN2[21] | select_n2x_1 & (~ IN2[21]) | select_ne_1 & (~ IN2[22])  );
    wire logic pp_1_23;
    assign pp_1_23 = (select_e_1 & IN2[23] | select_2x_1 & IN2[22] | select_n2x_1 & (~ IN2[22]) | select_ne_1 & (~ IN2[23])  );
    wire logic pp_1_24;
    assign pp_1_24 = (select_e_1 & IN2[24] | select_2x_1 & IN2[23] | select_n2x_1 & (~ IN2[23]) | select_ne_1 & (~ IN2[24])  );
    wire logic pp_1_25;
    assign pp_1_25 = (select_e_1 & IN2[25] | select_2x_1 & IN2[24] | select_n2x_1 & (~ IN2[24]) | select_ne_1 & (~ IN2[25])  );
    wire logic pp_1_26;
    assign pp_1_26 = (select_e_1 & IN2[26] | select_2x_1 & IN2[25] | select_n2x_1 & (~ IN2[25]) | select_ne_1 & (~ IN2[26])  );
    wire logic pp_1_27;
    assign pp_1_27 = (select_e_1 & IN2[27] | select_2x_1 & IN2[26] | select_n2x_1 & (~ IN2[26]) | select_ne_1 & (~ IN2[27])  );
    wire logic pp_1_28;
    assign pp_1_28 = (select_e_1 & IN2[28] | select_2x_1 & IN2[27] | select_n2x_1 & (~ IN2[27]) | select_ne_1 & (~ IN2[28])  );
    wire logic pp_1_29;
    assign pp_1_29 = (select_e_1 & IN2[29] | select_2x_1 & IN2[28] | select_n2x_1 & (~ IN2[28]) | select_ne_1 & (~ IN2[29])  );
    wire logic pp_1_30;
    assign pp_1_30 = (select_e_1 & IN2[30] | select_2x_1 & IN2[29] | select_n2x_1 & (~ IN2[29]) | select_ne_1 & (~ IN2[30])  );
    wire logic pp_1_31;
    assign pp_1_31 = (select_e_1 & IN2[31] | select_2x_1 & IN2[30] | select_n2x_1 & (~ IN2[30]) | select_ne_1 & (~ IN2[31])  );
    wire logic pp_1_32;
    assign pp_1_32 = (select_e_1 & IN2[32] | select_2x_1 & IN2[31] | select_n2x_1 & (~ IN2[31]) | select_ne_1 & (~ IN2[32])  );
    wire logic pp_1_33;
    assign pp_1_33 = (select_e_1 & IN2[33] | select_2x_1 & IN2[32] | select_n2x_1 & (~ IN2[32]) | select_ne_1 & (~ IN2[33])  );
    wire logic pp_1_34;
    assign pp_1_34 = (select_e_1 & IN2[34] | select_2x_1 & IN2[33] | select_n2x_1 & (~ IN2[33]) | select_ne_1 & (~ IN2[34])  );
    wire logic pp_1_35;
    assign pp_1_35 = (select_e_1 & IN2[35] | select_2x_1 & IN2[34] | select_n2x_1 & (~ IN2[34]) | select_ne_1 & (~ IN2[35])  );
    wire logic pp_1_36;
    assign pp_1_36 = (select_e_1 & IN2[36] | select_2x_1 & IN2[35] | select_n2x_1 & (~ IN2[35]) | select_ne_1 & (~ IN2[36])  );
    wire logic pp_1_37;
    assign pp_1_37 = (select_e_1 & IN2[37] | select_2x_1 & IN2[36] | select_n2x_1 & (~ IN2[36]) | select_ne_1 & (~ IN2[37])  );
    wire logic pp_1_38;
    assign pp_1_38 = (select_e_1 & IN2[38] | select_2x_1 & IN2[37] | select_n2x_1 & (~ IN2[37]) | select_ne_1 & (~ IN2[38])  );
    wire logic pp_1_39;
    assign pp_1_39 = (select_e_1 & IN2[39] | select_2x_1 & IN2[38] | select_n2x_1 & (~ IN2[38]) | select_ne_1 & (~ IN2[39])  );
    wire logic pp_1_40;
    assign pp_1_40 = (select_e_1 & IN2[40] | select_2x_1 & IN2[39] | select_n2x_1 & (~ IN2[39]) | select_ne_1 & (~ IN2[40])  );
    wire logic pp_1_41;
    assign pp_1_41 = (select_e_1 & IN2[41] | select_2x_1 & IN2[40] | select_n2x_1 & (~ IN2[40]) | select_ne_1 & (~ IN2[41])  );
    wire logic pp_1_42;
    assign pp_1_42 = (select_e_1 & IN2[42] | select_2x_1 & IN2[41] | select_n2x_1 & (~ IN2[41]) | select_ne_1 & (~ IN2[42])  );
    wire logic pp_1_43;
    assign pp_1_43 = (select_e_1 & IN2[43] | select_2x_1 & IN2[42] | select_n2x_1 & (~ IN2[42]) | select_ne_1 & (~ IN2[43])  );
    wire logic pp_1_44;
    assign pp_1_44 = (select_e_1 & IN2[44] | select_2x_1 & IN2[43] | select_n2x_1 & (~ IN2[43]) | select_ne_1 & (~ IN2[44])  );
    wire logic pp_1_45;
    assign pp_1_45 = (select_e_1 & IN2[45] | select_2x_1 & IN2[44] | select_n2x_1 & (~ IN2[44]) | select_ne_1 & (~ IN2[45])  );
    wire logic pp_1_46;
    assign pp_1_46 = (select_e_1 & IN2[46] | select_2x_1 & IN2[45] | select_n2x_1 & (~ IN2[45]) | select_ne_1 & (~ IN2[46])  );
    wire logic pp_1_47;
    assign pp_1_47 = (select_e_1 & IN2[47] | select_2x_1 & IN2[46] | select_n2x_1 & (~ IN2[46]) | select_ne_1 & (~ IN2[47])  );
    wire logic pp_1_48;
    assign pp_1_48 = (select_e_1 & IN2[48] | select_2x_1 & IN2[47] | select_n2x_1 & (~ IN2[47]) | select_ne_1 & (~ IN2[48])  );
    wire logic pp_1_49;
    assign pp_1_49 = (select_e_1 & IN2[49] | select_2x_1 & IN2[48] | select_n2x_1 & (~ IN2[48]) | select_ne_1 & (~ IN2[49])  );
    wire logic pp_1_50;
    assign pp_1_50 = (select_e_1 & IN2[50] | select_2x_1 & IN2[49] | select_n2x_1 & (~ IN2[49]) | select_ne_1 & (~ IN2[50])  );
    wire logic pp_1_51;
    assign pp_1_51 = (select_e_1 & IN2[51] | select_2x_1 & IN2[50] | select_n2x_1 & (~ IN2[50]) | select_ne_1 & (~ IN2[51])  );
    wire logic pp_1_52;
    assign pp_1_52 = (select_e_1 & IN2[52] | select_2x_1 & IN2[51] | select_n2x_1 & (~ IN2[51]) | select_ne_1 & (~ IN2[52])  );
    wire logic pp_1_53;
    assign pp_1_53 = (select_e_1 & IN2[53] | select_2x_1 & IN2[52] | select_n2x_1 & (~ IN2[52]) | select_ne_1 & (~ IN2[53])  );
    wire logic pp_1_54;
    assign pp_1_54 = (select_e_1 & IN2[54] | select_2x_1 & IN2[53] | select_n2x_1 & (~ IN2[53]) | select_ne_1 & (~ IN2[54])  );
    wire logic pp_1_55;
    assign pp_1_55 = (select_e_1 & IN2[55] | select_2x_1 & IN2[54] | select_n2x_1 & (~ IN2[54]) | select_ne_1 & (~ IN2[55])  );
    wire logic pp_1_56;
    assign pp_1_56 = (select_e_1 & IN2[56] | select_2x_1 & IN2[55] | select_n2x_1 & (~ IN2[55]) | select_ne_1 & (~ IN2[56])  );
    wire logic pp_1_57;
    assign pp_1_57 = (select_e_1 & IN2[57] | select_2x_1 & IN2[56] | select_n2x_1 & (~ IN2[56]) | select_ne_1 & (~ IN2[57])  );
    wire logic pp_1_58;
    assign pp_1_58 = (select_e_1 & IN2[58] | select_2x_1 & IN2[57] | select_n2x_1 & (~ IN2[57]) | select_ne_1 & (~ IN2[58])  );
    wire logic pp_1_59;
    assign pp_1_59 = (select_e_1 & IN2[59] | select_2x_1 & IN2[58] | select_n2x_1 & (~ IN2[58]) | select_ne_1 & (~ IN2[59])  );
    wire logic pp_1_60;
    assign pp_1_60 = (select_e_1 & IN2[60] | select_2x_1 & IN2[59] | select_n2x_1 & (~ IN2[59]) | select_ne_1 & (~ IN2[60])  );
    wire logic pp_1_61;
    assign pp_1_61 = (select_e_1 & IN2[61] | select_2x_1 & IN2[60] | select_n2x_1 & (~ IN2[60]) | select_ne_1 & (~ IN2[61])  );
    wire logic pp_1_62;
    assign pp_1_62 = (select_e_1 & IN2[62] | select_2x_1 & IN2[61] | select_n2x_1 & (~ IN2[61]) | select_ne_1 & (~ IN2[62])  );
    wire logic pp_1_63;
    assign pp_1_63 = (select_e_1 & IN2[63] | select_2x_1 & IN2[62] | select_n2x_1 & (~ IN2[62]) | select_ne_1 & (~ IN2[63])  );
    wire logic pp_1_64;
    assign pp_1_64 = (select_e_1 & IN2[63] | select_2x_1 & IN2[63] | select_n2x_1 & (~ IN2[63]) | select_ne_1 & (~ IN2[63])  );
    wire logic pp_1_65;
    assign pp_1_65 = ~ (select_e_1 & IN2[63] | select_2x_1 & IN2[63] | select_n2x_1 & (~ IN2[63]) | select_ne_1 & (~ IN2[63])  );
    assign tcomp1 = select_ne_1 | select_n2x_1;
    
    // Signed Booth Radix-4 Partial Products Row 3
    wire logic select_e_2, select_ne_2, select_2x_2, tcomp2, select_n2x_2;
    assign select_e_2 = ((~ IN1[5]) & (IN1[4] ^ IN1[3]));
    assign select_ne_2 = IN1[5] &  (IN1[4] ^ IN1[3]);
    assign select_2x_2 = (~ IN1[5]) & IN1[4] & IN1[3];
    assign select_n2x_2 = IN1[5] & (~ IN1[4]) & (~ IN1[3]);
    wire logic pp_2_0;
    assign pp_2_0 = (select_e_2 & IN2[0] | select_2x_2 & 1'b0 | select_n2x_2 & 1'b1 | select_ne_2 & (~ IN2[0])  );
    wire logic pp_2_1;
    assign pp_2_1 = (select_e_2 & IN2[1] | select_2x_2 & IN2[0] | select_n2x_2 & (~ IN2[0]) | select_ne_2 & (~ IN2[1])  );
    wire logic pp_2_2;
    assign pp_2_2 = (select_e_2 & IN2[2] | select_2x_2 & IN2[1] | select_n2x_2 & (~ IN2[1]) | select_ne_2 & (~ IN2[2])  );
    wire logic pp_2_3;
    assign pp_2_3 = (select_e_2 & IN2[3] | select_2x_2 & IN2[2] | select_n2x_2 & (~ IN2[2]) | select_ne_2 & (~ IN2[3])  );
    wire logic pp_2_4;
    assign pp_2_4 = (select_e_2 & IN2[4] | select_2x_2 & IN2[3] | select_n2x_2 & (~ IN2[3]) | select_ne_2 & (~ IN2[4])  );
    wire logic pp_2_5;
    assign pp_2_5 = (select_e_2 & IN2[5] | select_2x_2 & IN2[4] | select_n2x_2 & (~ IN2[4]) | select_ne_2 & (~ IN2[5])  );
    wire logic pp_2_6;
    assign pp_2_6 = (select_e_2 & IN2[6] | select_2x_2 & IN2[5] | select_n2x_2 & (~ IN2[5]) | select_ne_2 & (~ IN2[6])  );
    wire logic pp_2_7;
    assign pp_2_7 = (select_e_2 & IN2[7] | select_2x_2 & IN2[6] | select_n2x_2 & (~ IN2[6]) | select_ne_2 & (~ IN2[7])  );
    wire logic pp_2_8;
    assign pp_2_8 = (select_e_2 & IN2[8] | select_2x_2 & IN2[7] | select_n2x_2 & (~ IN2[7]) | select_ne_2 & (~ IN2[8])  );
    wire logic pp_2_9;
    assign pp_2_9 = (select_e_2 & IN2[9] | select_2x_2 & IN2[8] | select_n2x_2 & (~ IN2[8]) | select_ne_2 & (~ IN2[9])  );
    wire logic pp_2_10;
    assign pp_2_10 = (select_e_2 & IN2[10] | select_2x_2 & IN2[9] | select_n2x_2 & (~ IN2[9]) | select_ne_2 & (~ IN2[10])  );
    wire logic pp_2_11;
    assign pp_2_11 = (select_e_2 & IN2[11] | select_2x_2 & IN2[10] | select_n2x_2 & (~ IN2[10]) | select_ne_2 & (~ IN2[11])  );
    wire logic pp_2_12;
    assign pp_2_12 = (select_e_2 & IN2[12] | select_2x_2 & IN2[11] | select_n2x_2 & (~ IN2[11]) | select_ne_2 & (~ IN2[12])  );
    wire logic pp_2_13;
    assign pp_2_13 = (select_e_2 & IN2[13] | select_2x_2 & IN2[12] | select_n2x_2 & (~ IN2[12]) | select_ne_2 & (~ IN2[13])  );
    wire logic pp_2_14;
    assign pp_2_14 = (select_e_2 & IN2[14] | select_2x_2 & IN2[13] | select_n2x_2 & (~ IN2[13]) | select_ne_2 & (~ IN2[14])  );
    wire logic pp_2_15;
    assign pp_2_15 = (select_e_2 & IN2[15] | select_2x_2 & IN2[14] | select_n2x_2 & (~ IN2[14]) | select_ne_2 & (~ IN2[15])  );
    wire logic pp_2_16;
    assign pp_2_16 = (select_e_2 & IN2[16] | select_2x_2 & IN2[15] | select_n2x_2 & (~ IN2[15]) | select_ne_2 & (~ IN2[16])  );
    wire logic pp_2_17;
    assign pp_2_17 = (select_e_2 & IN2[17] | select_2x_2 & IN2[16] | select_n2x_2 & (~ IN2[16]) | select_ne_2 & (~ IN2[17])  );
    wire logic pp_2_18;
    assign pp_2_18 = (select_e_2 & IN2[18] | select_2x_2 & IN2[17] | select_n2x_2 & (~ IN2[17]) | select_ne_2 & (~ IN2[18])  );
    wire logic pp_2_19;
    assign pp_2_19 = (select_e_2 & IN2[19] | select_2x_2 & IN2[18] | select_n2x_2 & (~ IN2[18]) | select_ne_2 & (~ IN2[19])  );
    wire logic pp_2_20;
    assign pp_2_20 = (select_e_2 & IN2[20] | select_2x_2 & IN2[19] | select_n2x_2 & (~ IN2[19]) | select_ne_2 & (~ IN2[20])  );
    wire logic pp_2_21;
    assign pp_2_21 = (select_e_2 & IN2[21] | select_2x_2 & IN2[20] | select_n2x_2 & (~ IN2[20]) | select_ne_2 & (~ IN2[21])  );
    wire logic pp_2_22;
    assign pp_2_22 = (select_e_2 & IN2[22] | select_2x_2 & IN2[21] | select_n2x_2 & (~ IN2[21]) | select_ne_2 & (~ IN2[22])  );
    wire logic pp_2_23;
    assign pp_2_23 = (select_e_2 & IN2[23] | select_2x_2 & IN2[22] | select_n2x_2 & (~ IN2[22]) | select_ne_2 & (~ IN2[23])  );
    wire logic pp_2_24;
    assign pp_2_24 = (select_e_2 & IN2[24] | select_2x_2 & IN2[23] | select_n2x_2 & (~ IN2[23]) | select_ne_2 & (~ IN2[24])  );
    wire logic pp_2_25;
    assign pp_2_25 = (select_e_2 & IN2[25] | select_2x_2 & IN2[24] | select_n2x_2 & (~ IN2[24]) | select_ne_2 & (~ IN2[25])  );
    wire logic pp_2_26;
    assign pp_2_26 = (select_e_2 & IN2[26] | select_2x_2 & IN2[25] | select_n2x_2 & (~ IN2[25]) | select_ne_2 & (~ IN2[26])  );
    wire logic pp_2_27;
    assign pp_2_27 = (select_e_2 & IN2[27] | select_2x_2 & IN2[26] | select_n2x_2 & (~ IN2[26]) | select_ne_2 & (~ IN2[27])  );
    wire logic pp_2_28;
    assign pp_2_28 = (select_e_2 & IN2[28] | select_2x_2 & IN2[27] | select_n2x_2 & (~ IN2[27]) | select_ne_2 & (~ IN2[28])  );
    wire logic pp_2_29;
    assign pp_2_29 = (select_e_2 & IN2[29] | select_2x_2 & IN2[28] | select_n2x_2 & (~ IN2[28]) | select_ne_2 & (~ IN2[29])  );
    wire logic pp_2_30;
    assign pp_2_30 = (select_e_2 & IN2[30] | select_2x_2 & IN2[29] | select_n2x_2 & (~ IN2[29]) | select_ne_2 & (~ IN2[30])  );
    wire logic pp_2_31;
    assign pp_2_31 = (select_e_2 & IN2[31] | select_2x_2 & IN2[30] | select_n2x_2 & (~ IN2[30]) | select_ne_2 & (~ IN2[31])  );
    wire logic pp_2_32;
    assign pp_2_32 = (select_e_2 & IN2[32] | select_2x_2 & IN2[31] | select_n2x_2 & (~ IN2[31]) | select_ne_2 & (~ IN2[32])  );
    wire logic pp_2_33;
    assign pp_2_33 = (select_e_2 & IN2[33] | select_2x_2 & IN2[32] | select_n2x_2 & (~ IN2[32]) | select_ne_2 & (~ IN2[33])  );
    wire logic pp_2_34;
    assign pp_2_34 = (select_e_2 & IN2[34] | select_2x_2 & IN2[33] | select_n2x_2 & (~ IN2[33]) | select_ne_2 & (~ IN2[34])  );
    wire logic pp_2_35;
    assign pp_2_35 = (select_e_2 & IN2[35] | select_2x_2 & IN2[34] | select_n2x_2 & (~ IN2[34]) | select_ne_2 & (~ IN2[35])  );
    wire logic pp_2_36;
    assign pp_2_36 = (select_e_2 & IN2[36] | select_2x_2 & IN2[35] | select_n2x_2 & (~ IN2[35]) | select_ne_2 & (~ IN2[36])  );
    wire logic pp_2_37;
    assign pp_2_37 = (select_e_2 & IN2[37] | select_2x_2 & IN2[36] | select_n2x_2 & (~ IN2[36]) | select_ne_2 & (~ IN2[37])  );
    wire logic pp_2_38;
    assign pp_2_38 = (select_e_2 & IN2[38] | select_2x_2 & IN2[37] | select_n2x_2 & (~ IN2[37]) | select_ne_2 & (~ IN2[38])  );
    wire logic pp_2_39;
    assign pp_2_39 = (select_e_2 & IN2[39] | select_2x_2 & IN2[38] | select_n2x_2 & (~ IN2[38]) | select_ne_2 & (~ IN2[39])  );
    wire logic pp_2_40;
    assign pp_2_40 = (select_e_2 & IN2[40] | select_2x_2 & IN2[39] | select_n2x_2 & (~ IN2[39]) | select_ne_2 & (~ IN2[40])  );
    wire logic pp_2_41;
    assign pp_2_41 = (select_e_2 & IN2[41] | select_2x_2 & IN2[40] | select_n2x_2 & (~ IN2[40]) | select_ne_2 & (~ IN2[41])  );
    wire logic pp_2_42;
    assign pp_2_42 = (select_e_2 & IN2[42] | select_2x_2 & IN2[41] | select_n2x_2 & (~ IN2[41]) | select_ne_2 & (~ IN2[42])  );
    wire logic pp_2_43;
    assign pp_2_43 = (select_e_2 & IN2[43] | select_2x_2 & IN2[42] | select_n2x_2 & (~ IN2[42]) | select_ne_2 & (~ IN2[43])  );
    wire logic pp_2_44;
    assign pp_2_44 = (select_e_2 & IN2[44] | select_2x_2 & IN2[43] | select_n2x_2 & (~ IN2[43]) | select_ne_2 & (~ IN2[44])  );
    wire logic pp_2_45;
    assign pp_2_45 = (select_e_2 & IN2[45] | select_2x_2 & IN2[44] | select_n2x_2 & (~ IN2[44]) | select_ne_2 & (~ IN2[45])  );
    wire logic pp_2_46;
    assign pp_2_46 = (select_e_2 & IN2[46] | select_2x_2 & IN2[45] | select_n2x_2 & (~ IN2[45]) | select_ne_2 & (~ IN2[46])  );
    wire logic pp_2_47;
    assign pp_2_47 = (select_e_2 & IN2[47] | select_2x_2 & IN2[46] | select_n2x_2 & (~ IN2[46]) | select_ne_2 & (~ IN2[47])  );
    wire logic pp_2_48;
    assign pp_2_48 = (select_e_2 & IN2[48] | select_2x_2 & IN2[47] | select_n2x_2 & (~ IN2[47]) | select_ne_2 & (~ IN2[48])  );
    wire logic pp_2_49;
    assign pp_2_49 = (select_e_2 & IN2[49] | select_2x_2 & IN2[48] | select_n2x_2 & (~ IN2[48]) | select_ne_2 & (~ IN2[49])  );
    wire logic pp_2_50;
    assign pp_2_50 = (select_e_2 & IN2[50] | select_2x_2 & IN2[49] | select_n2x_2 & (~ IN2[49]) | select_ne_2 & (~ IN2[50])  );
    wire logic pp_2_51;
    assign pp_2_51 = (select_e_2 & IN2[51] | select_2x_2 & IN2[50] | select_n2x_2 & (~ IN2[50]) | select_ne_2 & (~ IN2[51])  );
    wire logic pp_2_52;
    assign pp_2_52 = (select_e_2 & IN2[52] | select_2x_2 & IN2[51] | select_n2x_2 & (~ IN2[51]) | select_ne_2 & (~ IN2[52])  );
    wire logic pp_2_53;
    assign pp_2_53 = (select_e_2 & IN2[53] | select_2x_2 & IN2[52] | select_n2x_2 & (~ IN2[52]) | select_ne_2 & (~ IN2[53])  );
    wire logic pp_2_54;
    assign pp_2_54 = (select_e_2 & IN2[54] | select_2x_2 & IN2[53] | select_n2x_2 & (~ IN2[53]) | select_ne_2 & (~ IN2[54])  );
    wire logic pp_2_55;
    assign pp_2_55 = (select_e_2 & IN2[55] | select_2x_2 & IN2[54] | select_n2x_2 & (~ IN2[54]) | select_ne_2 & (~ IN2[55])  );
    wire logic pp_2_56;
    assign pp_2_56 = (select_e_2 & IN2[56] | select_2x_2 & IN2[55] | select_n2x_2 & (~ IN2[55]) | select_ne_2 & (~ IN2[56])  );
    wire logic pp_2_57;
    assign pp_2_57 = (select_e_2 & IN2[57] | select_2x_2 & IN2[56] | select_n2x_2 & (~ IN2[56]) | select_ne_2 & (~ IN2[57])  );
    wire logic pp_2_58;
    assign pp_2_58 = (select_e_2 & IN2[58] | select_2x_2 & IN2[57] | select_n2x_2 & (~ IN2[57]) | select_ne_2 & (~ IN2[58])  );
    wire logic pp_2_59;
    assign pp_2_59 = (select_e_2 & IN2[59] | select_2x_2 & IN2[58] | select_n2x_2 & (~ IN2[58]) | select_ne_2 & (~ IN2[59])  );
    wire logic pp_2_60;
    assign pp_2_60 = (select_e_2 & IN2[60] | select_2x_2 & IN2[59] | select_n2x_2 & (~ IN2[59]) | select_ne_2 & (~ IN2[60])  );
    wire logic pp_2_61;
    assign pp_2_61 = (select_e_2 & IN2[61] | select_2x_2 & IN2[60] | select_n2x_2 & (~ IN2[60]) | select_ne_2 & (~ IN2[61])  );
    wire logic pp_2_62;
    assign pp_2_62 = (select_e_2 & IN2[62] | select_2x_2 & IN2[61] | select_n2x_2 & (~ IN2[61]) | select_ne_2 & (~ IN2[62])  );
    wire logic pp_2_63;
    assign pp_2_63 = (select_e_2 & IN2[63] | select_2x_2 & IN2[62] | select_n2x_2 & (~ IN2[62]) | select_ne_2 & (~ IN2[63])  );
    wire logic pp_2_64;
    assign pp_2_64 = (select_e_2 & IN2[63] | select_2x_2 & IN2[63] | select_n2x_2 & (~ IN2[63]) | select_ne_2 & (~ IN2[63])  );
    wire logic pp_2_65;
    assign pp_2_65 = ~ (select_e_2 & IN2[63] | select_2x_2 & IN2[63] | select_n2x_2 & (~ IN2[63]) | select_ne_2 & (~ IN2[63])  );
    assign tcomp2 = select_ne_2 | select_n2x_2;
    
    // Signed Booth Radix-4 Partial Products Row 4
    wire logic select_e_3, select_ne_3, select_2x_3, tcomp3, select_n2x_3;
    assign select_e_3 = ((~ IN1[7]) & (IN1[6] ^ IN1[5]));
    assign select_ne_3 = IN1[7] &  (IN1[6] ^ IN1[5]);
    assign select_2x_3 = (~ IN1[7]) & IN1[6] & IN1[5];
    assign select_n2x_3 = IN1[7] & (~ IN1[6]) & (~ IN1[5]);
    wire logic pp_3_0;
    assign pp_3_0 = (select_e_3 & IN2[0] | select_2x_3 & 1'b0 | select_n2x_3 & 1'b1 | select_ne_3 & (~ IN2[0])  );
    wire logic pp_3_1;
    assign pp_3_1 = (select_e_3 & IN2[1] | select_2x_3 & IN2[0] | select_n2x_3 & (~ IN2[0]) | select_ne_3 & (~ IN2[1])  );
    wire logic pp_3_2;
    assign pp_3_2 = (select_e_3 & IN2[2] | select_2x_3 & IN2[1] | select_n2x_3 & (~ IN2[1]) | select_ne_3 & (~ IN2[2])  );
    wire logic pp_3_3;
    assign pp_3_3 = (select_e_3 & IN2[3] | select_2x_3 & IN2[2] | select_n2x_3 & (~ IN2[2]) | select_ne_3 & (~ IN2[3])  );
    wire logic pp_3_4;
    assign pp_3_4 = (select_e_3 & IN2[4] | select_2x_3 & IN2[3] | select_n2x_3 & (~ IN2[3]) | select_ne_3 & (~ IN2[4])  );
    wire logic pp_3_5;
    assign pp_3_5 = (select_e_3 & IN2[5] | select_2x_3 & IN2[4] | select_n2x_3 & (~ IN2[4]) | select_ne_3 & (~ IN2[5])  );
    wire logic pp_3_6;
    assign pp_3_6 = (select_e_3 & IN2[6] | select_2x_3 & IN2[5] | select_n2x_3 & (~ IN2[5]) | select_ne_3 & (~ IN2[6])  );
    wire logic pp_3_7;
    assign pp_3_7 = (select_e_3 & IN2[7] | select_2x_3 & IN2[6] | select_n2x_3 & (~ IN2[6]) | select_ne_3 & (~ IN2[7])  );
    wire logic pp_3_8;
    assign pp_3_8 = (select_e_3 & IN2[8] | select_2x_3 & IN2[7] | select_n2x_3 & (~ IN2[7]) | select_ne_3 & (~ IN2[8])  );
    wire logic pp_3_9;
    assign pp_3_9 = (select_e_3 & IN2[9] | select_2x_3 & IN2[8] | select_n2x_3 & (~ IN2[8]) | select_ne_3 & (~ IN2[9])  );
    wire logic pp_3_10;
    assign pp_3_10 = (select_e_3 & IN2[10] | select_2x_3 & IN2[9] | select_n2x_3 & (~ IN2[9]) | select_ne_3 & (~ IN2[10])  );
    wire logic pp_3_11;
    assign pp_3_11 = (select_e_3 & IN2[11] | select_2x_3 & IN2[10] | select_n2x_3 & (~ IN2[10]) | select_ne_3 & (~ IN2[11])  );
    wire logic pp_3_12;
    assign pp_3_12 = (select_e_3 & IN2[12] | select_2x_3 & IN2[11] | select_n2x_3 & (~ IN2[11]) | select_ne_3 & (~ IN2[12])  );
    wire logic pp_3_13;
    assign pp_3_13 = (select_e_3 & IN2[13] | select_2x_3 & IN2[12] | select_n2x_3 & (~ IN2[12]) | select_ne_3 & (~ IN2[13])  );
    wire logic pp_3_14;
    assign pp_3_14 = (select_e_3 & IN2[14] | select_2x_3 & IN2[13] | select_n2x_3 & (~ IN2[13]) | select_ne_3 & (~ IN2[14])  );
    wire logic pp_3_15;
    assign pp_3_15 = (select_e_3 & IN2[15] | select_2x_3 & IN2[14] | select_n2x_3 & (~ IN2[14]) | select_ne_3 & (~ IN2[15])  );
    wire logic pp_3_16;
    assign pp_3_16 = (select_e_3 & IN2[16] | select_2x_3 & IN2[15] | select_n2x_3 & (~ IN2[15]) | select_ne_3 & (~ IN2[16])  );
    wire logic pp_3_17;
    assign pp_3_17 = (select_e_3 & IN2[17] | select_2x_3 & IN2[16] | select_n2x_3 & (~ IN2[16]) | select_ne_3 & (~ IN2[17])  );
    wire logic pp_3_18;
    assign pp_3_18 = (select_e_3 & IN2[18] | select_2x_3 & IN2[17] | select_n2x_3 & (~ IN2[17]) | select_ne_3 & (~ IN2[18])  );
    wire logic pp_3_19;
    assign pp_3_19 = (select_e_3 & IN2[19] | select_2x_3 & IN2[18] | select_n2x_3 & (~ IN2[18]) | select_ne_3 & (~ IN2[19])  );
    wire logic pp_3_20;
    assign pp_3_20 = (select_e_3 & IN2[20] | select_2x_3 & IN2[19] | select_n2x_3 & (~ IN2[19]) | select_ne_3 & (~ IN2[20])  );
    wire logic pp_3_21;
    assign pp_3_21 = (select_e_3 & IN2[21] | select_2x_3 & IN2[20] | select_n2x_3 & (~ IN2[20]) | select_ne_3 & (~ IN2[21])  );
    wire logic pp_3_22;
    assign pp_3_22 = (select_e_3 & IN2[22] | select_2x_3 & IN2[21] | select_n2x_3 & (~ IN2[21]) | select_ne_3 & (~ IN2[22])  );
    wire logic pp_3_23;
    assign pp_3_23 = (select_e_3 & IN2[23] | select_2x_3 & IN2[22] | select_n2x_3 & (~ IN2[22]) | select_ne_3 & (~ IN2[23])  );
    wire logic pp_3_24;
    assign pp_3_24 = (select_e_3 & IN2[24] | select_2x_3 & IN2[23] | select_n2x_3 & (~ IN2[23]) | select_ne_3 & (~ IN2[24])  );
    wire logic pp_3_25;
    assign pp_3_25 = (select_e_3 & IN2[25] | select_2x_3 & IN2[24] | select_n2x_3 & (~ IN2[24]) | select_ne_3 & (~ IN2[25])  );
    wire logic pp_3_26;
    assign pp_3_26 = (select_e_3 & IN2[26] | select_2x_3 & IN2[25] | select_n2x_3 & (~ IN2[25]) | select_ne_3 & (~ IN2[26])  );
    wire logic pp_3_27;
    assign pp_3_27 = (select_e_3 & IN2[27] | select_2x_3 & IN2[26] | select_n2x_3 & (~ IN2[26]) | select_ne_3 & (~ IN2[27])  );
    wire logic pp_3_28;
    assign pp_3_28 = (select_e_3 & IN2[28] | select_2x_3 & IN2[27] | select_n2x_3 & (~ IN2[27]) | select_ne_3 & (~ IN2[28])  );
    wire logic pp_3_29;
    assign pp_3_29 = (select_e_3 & IN2[29] | select_2x_3 & IN2[28] | select_n2x_3 & (~ IN2[28]) | select_ne_3 & (~ IN2[29])  );
    wire logic pp_3_30;
    assign pp_3_30 = (select_e_3 & IN2[30] | select_2x_3 & IN2[29] | select_n2x_3 & (~ IN2[29]) | select_ne_3 & (~ IN2[30])  );
    wire logic pp_3_31;
    assign pp_3_31 = (select_e_3 & IN2[31] | select_2x_3 & IN2[30] | select_n2x_3 & (~ IN2[30]) | select_ne_3 & (~ IN2[31])  );
    wire logic pp_3_32;
    assign pp_3_32 = (select_e_3 & IN2[32] | select_2x_3 & IN2[31] | select_n2x_3 & (~ IN2[31]) | select_ne_3 & (~ IN2[32])  );
    wire logic pp_3_33;
    assign pp_3_33 = (select_e_3 & IN2[33] | select_2x_3 & IN2[32] | select_n2x_3 & (~ IN2[32]) | select_ne_3 & (~ IN2[33])  );
    wire logic pp_3_34;
    assign pp_3_34 = (select_e_3 & IN2[34] | select_2x_3 & IN2[33] | select_n2x_3 & (~ IN2[33]) | select_ne_3 & (~ IN2[34])  );
    wire logic pp_3_35;
    assign pp_3_35 = (select_e_3 & IN2[35] | select_2x_3 & IN2[34] | select_n2x_3 & (~ IN2[34]) | select_ne_3 & (~ IN2[35])  );
    wire logic pp_3_36;
    assign pp_3_36 = (select_e_3 & IN2[36] | select_2x_3 & IN2[35] | select_n2x_3 & (~ IN2[35]) | select_ne_3 & (~ IN2[36])  );
    wire logic pp_3_37;
    assign pp_3_37 = (select_e_3 & IN2[37] | select_2x_3 & IN2[36] | select_n2x_3 & (~ IN2[36]) | select_ne_3 & (~ IN2[37])  );
    wire logic pp_3_38;
    assign pp_3_38 = (select_e_3 & IN2[38] | select_2x_3 & IN2[37] | select_n2x_3 & (~ IN2[37]) | select_ne_3 & (~ IN2[38])  );
    wire logic pp_3_39;
    assign pp_3_39 = (select_e_3 & IN2[39] | select_2x_3 & IN2[38] | select_n2x_3 & (~ IN2[38]) | select_ne_3 & (~ IN2[39])  );
    wire logic pp_3_40;
    assign pp_3_40 = (select_e_3 & IN2[40] | select_2x_3 & IN2[39] | select_n2x_3 & (~ IN2[39]) | select_ne_3 & (~ IN2[40])  );
    wire logic pp_3_41;
    assign pp_3_41 = (select_e_3 & IN2[41] | select_2x_3 & IN2[40] | select_n2x_3 & (~ IN2[40]) | select_ne_3 & (~ IN2[41])  );
    wire logic pp_3_42;
    assign pp_3_42 = (select_e_3 & IN2[42] | select_2x_3 & IN2[41] | select_n2x_3 & (~ IN2[41]) | select_ne_3 & (~ IN2[42])  );
    wire logic pp_3_43;
    assign pp_3_43 = (select_e_3 & IN2[43] | select_2x_3 & IN2[42] | select_n2x_3 & (~ IN2[42]) | select_ne_3 & (~ IN2[43])  );
    wire logic pp_3_44;
    assign pp_3_44 = (select_e_3 & IN2[44] | select_2x_3 & IN2[43] | select_n2x_3 & (~ IN2[43]) | select_ne_3 & (~ IN2[44])  );
    wire logic pp_3_45;
    assign pp_3_45 = (select_e_3 & IN2[45] | select_2x_3 & IN2[44] | select_n2x_3 & (~ IN2[44]) | select_ne_3 & (~ IN2[45])  );
    wire logic pp_3_46;
    assign pp_3_46 = (select_e_3 & IN2[46] | select_2x_3 & IN2[45] | select_n2x_3 & (~ IN2[45]) | select_ne_3 & (~ IN2[46])  );
    wire logic pp_3_47;
    assign pp_3_47 = (select_e_3 & IN2[47] | select_2x_3 & IN2[46] | select_n2x_3 & (~ IN2[46]) | select_ne_3 & (~ IN2[47])  );
    wire logic pp_3_48;
    assign pp_3_48 = (select_e_3 & IN2[48] | select_2x_3 & IN2[47] | select_n2x_3 & (~ IN2[47]) | select_ne_3 & (~ IN2[48])  );
    wire logic pp_3_49;
    assign pp_3_49 = (select_e_3 & IN2[49] | select_2x_3 & IN2[48] | select_n2x_3 & (~ IN2[48]) | select_ne_3 & (~ IN2[49])  );
    wire logic pp_3_50;
    assign pp_3_50 = (select_e_3 & IN2[50] | select_2x_3 & IN2[49] | select_n2x_3 & (~ IN2[49]) | select_ne_3 & (~ IN2[50])  );
    wire logic pp_3_51;
    assign pp_3_51 = (select_e_3 & IN2[51] | select_2x_3 & IN2[50] | select_n2x_3 & (~ IN2[50]) | select_ne_3 & (~ IN2[51])  );
    wire logic pp_3_52;
    assign pp_3_52 = (select_e_3 & IN2[52] | select_2x_3 & IN2[51] | select_n2x_3 & (~ IN2[51]) | select_ne_3 & (~ IN2[52])  );
    wire logic pp_3_53;
    assign pp_3_53 = (select_e_3 & IN2[53] | select_2x_3 & IN2[52] | select_n2x_3 & (~ IN2[52]) | select_ne_3 & (~ IN2[53])  );
    wire logic pp_3_54;
    assign pp_3_54 = (select_e_3 & IN2[54] | select_2x_3 & IN2[53] | select_n2x_3 & (~ IN2[53]) | select_ne_3 & (~ IN2[54])  );
    wire logic pp_3_55;
    assign pp_3_55 = (select_e_3 & IN2[55] | select_2x_3 & IN2[54] | select_n2x_3 & (~ IN2[54]) | select_ne_3 & (~ IN2[55])  );
    wire logic pp_3_56;
    assign pp_3_56 = (select_e_3 & IN2[56] | select_2x_3 & IN2[55] | select_n2x_3 & (~ IN2[55]) | select_ne_3 & (~ IN2[56])  );
    wire logic pp_3_57;
    assign pp_3_57 = (select_e_3 & IN2[57] | select_2x_3 & IN2[56] | select_n2x_3 & (~ IN2[56]) | select_ne_3 & (~ IN2[57])  );
    wire logic pp_3_58;
    assign pp_3_58 = (select_e_3 & IN2[58] | select_2x_3 & IN2[57] | select_n2x_3 & (~ IN2[57]) | select_ne_3 & (~ IN2[58])  );
    wire logic pp_3_59;
    assign pp_3_59 = (select_e_3 & IN2[59] | select_2x_3 & IN2[58] | select_n2x_3 & (~ IN2[58]) | select_ne_3 & (~ IN2[59])  );
    wire logic pp_3_60;
    assign pp_3_60 = (select_e_3 & IN2[60] | select_2x_3 & IN2[59] | select_n2x_3 & (~ IN2[59]) | select_ne_3 & (~ IN2[60])  );
    wire logic pp_3_61;
    assign pp_3_61 = (select_e_3 & IN2[61] | select_2x_3 & IN2[60] | select_n2x_3 & (~ IN2[60]) | select_ne_3 & (~ IN2[61])  );
    wire logic pp_3_62;
    assign pp_3_62 = (select_e_3 & IN2[62] | select_2x_3 & IN2[61] | select_n2x_3 & (~ IN2[61]) | select_ne_3 & (~ IN2[62])  );
    wire logic pp_3_63;
    assign pp_3_63 = (select_e_3 & IN2[63] | select_2x_3 & IN2[62] | select_n2x_3 & (~ IN2[62]) | select_ne_3 & (~ IN2[63])  );
    wire logic pp_3_64;
    assign pp_3_64 = (select_e_3 & IN2[63] | select_2x_3 & IN2[63] | select_n2x_3 & (~ IN2[63]) | select_ne_3 & (~ IN2[63])  );
    wire logic pp_3_65;
    assign pp_3_65 = ~ (select_e_3 & IN2[63] | select_2x_3 & IN2[63] | select_n2x_3 & (~ IN2[63]) | select_ne_3 & (~ IN2[63])  );
    assign tcomp3 = select_ne_3 | select_n2x_3;
    
    // Signed Booth Radix-4 Partial Products Row 5
    wire logic select_e_4, select_ne_4, select_2x_4, tcomp4, select_n2x_4;
    assign select_e_4 = ((~ IN1[9]) & (IN1[8] ^ IN1[7]));
    assign select_ne_4 = IN1[9] &  (IN1[8] ^ IN1[7]);
    assign select_2x_4 = (~ IN1[9]) & IN1[8] & IN1[7];
    assign select_n2x_4 = IN1[9] & (~ IN1[8]) & (~ IN1[7]);
    wire logic pp_4_0;
    assign pp_4_0 = (select_e_4 & IN2[0] | select_2x_4 & 1'b0 | select_n2x_4 & 1'b1 | select_ne_4 & (~ IN2[0])  );
    wire logic pp_4_1;
    assign pp_4_1 = (select_e_4 & IN2[1] | select_2x_4 & IN2[0] | select_n2x_4 & (~ IN2[0]) | select_ne_4 & (~ IN2[1])  );
    wire logic pp_4_2;
    assign pp_4_2 = (select_e_4 & IN2[2] | select_2x_4 & IN2[1] | select_n2x_4 & (~ IN2[1]) | select_ne_4 & (~ IN2[2])  );
    wire logic pp_4_3;
    assign pp_4_3 = (select_e_4 & IN2[3] | select_2x_4 & IN2[2] | select_n2x_4 & (~ IN2[2]) | select_ne_4 & (~ IN2[3])  );
    wire logic pp_4_4;
    assign pp_4_4 = (select_e_4 & IN2[4] | select_2x_4 & IN2[3] | select_n2x_4 & (~ IN2[3]) | select_ne_4 & (~ IN2[4])  );
    wire logic pp_4_5;
    assign pp_4_5 = (select_e_4 & IN2[5] | select_2x_4 & IN2[4] | select_n2x_4 & (~ IN2[4]) | select_ne_4 & (~ IN2[5])  );
    wire logic pp_4_6;
    assign pp_4_6 = (select_e_4 & IN2[6] | select_2x_4 & IN2[5] | select_n2x_4 & (~ IN2[5]) | select_ne_4 & (~ IN2[6])  );
    wire logic pp_4_7;
    assign pp_4_7 = (select_e_4 & IN2[7] | select_2x_4 & IN2[6] | select_n2x_4 & (~ IN2[6]) | select_ne_4 & (~ IN2[7])  );
    wire logic pp_4_8;
    assign pp_4_8 = (select_e_4 & IN2[8] | select_2x_4 & IN2[7] | select_n2x_4 & (~ IN2[7]) | select_ne_4 & (~ IN2[8])  );
    wire logic pp_4_9;
    assign pp_4_9 = (select_e_4 & IN2[9] | select_2x_4 & IN2[8] | select_n2x_4 & (~ IN2[8]) | select_ne_4 & (~ IN2[9])  );
    wire logic pp_4_10;
    assign pp_4_10 = (select_e_4 & IN2[10] | select_2x_4 & IN2[9] | select_n2x_4 & (~ IN2[9]) | select_ne_4 & (~ IN2[10])  );
    wire logic pp_4_11;
    assign pp_4_11 = (select_e_4 & IN2[11] | select_2x_4 & IN2[10] | select_n2x_4 & (~ IN2[10]) | select_ne_4 & (~ IN2[11])  );
    wire logic pp_4_12;
    assign pp_4_12 = (select_e_4 & IN2[12] | select_2x_4 & IN2[11] | select_n2x_4 & (~ IN2[11]) | select_ne_4 & (~ IN2[12])  );
    wire logic pp_4_13;
    assign pp_4_13 = (select_e_4 & IN2[13] | select_2x_4 & IN2[12] | select_n2x_4 & (~ IN2[12]) | select_ne_4 & (~ IN2[13])  );
    wire logic pp_4_14;
    assign pp_4_14 = (select_e_4 & IN2[14] | select_2x_4 & IN2[13] | select_n2x_4 & (~ IN2[13]) | select_ne_4 & (~ IN2[14])  );
    wire logic pp_4_15;
    assign pp_4_15 = (select_e_4 & IN2[15] | select_2x_4 & IN2[14] | select_n2x_4 & (~ IN2[14]) | select_ne_4 & (~ IN2[15])  );
    wire logic pp_4_16;
    assign pp_4_16 = (select_e_4 & IN2[16] | select_2x_4 & IN2[15] | select_n2x_4 & (~ IN2[15]) | select_ne_4 & (~ IN2[16])  );
    wire logic pp_4_17;
    assign pp_4_17 = (select_e_4 & IN2[17] | select_2x_4 & IN2[16] | select_n2x_4 & (~ IN2[16]) | select_ne_4 & (~ IN2[17])  );
    wire logic pp_4_18;
    assign pp_4_18 = (select_e_4 & IN2[18] | select_2x_4 & IN2[17] | select_n2x_4 & (~ IN2[17]) | select_ne_4 & (~ IN2[18])  );
    wire logic pp_4_19;
    assign pp_4_19 = (select_e_4 & IN2[19] | select_2x_4 & IN2[18] | select_n2x_4 & (~ IN2[18]) | select_ne_4 & (~ IN2[19])  );
    wire logic pp_4_20;
    assign pp_4_20 = (select_e_4 & IN2[20] | select_2x_4 & IN2[19] | select_n2x_4 & (~ IN2[19]) | select_ne_4 & (~ IN2[20])  );
    wire logic pp_4_21;
    assign pp_4_21 = (select_e_4 & IN2[21] | select_2x_4 & IN2[20] | select_n2x_4 & (~ IN2[20]) | select_ne_4 & (~ IN2[21])  );
    wire logic pp_4_22;
    assign pp_4_22 = (select_e_4 & IN2[22] | select_2x_4 & IN2[21] | select_n2x_4 & (~ IN2[21]) | select_ne_4 & (~ IN2[22])  );
    wire logic pp_4_23;
    assign pp_4_23 = (select_e_4 & IN2[23] | select_2x_4 & IN2[22] | select_n2x_4 & (~ IN2[22]) | select_ne_4 & (~ IN2[23])  );
    wire logic pp_4_24;
    assign pp_4_24 = (select_e_4 & IN2[24] | select_2x_4 & IN2[23] | select_n2x_4 & (~ IN2[23]) | select_ne_4 & (~ IN2[24])  );
    wire logic pp_4_25;
    assign pp_4_25 = (select_e_4 & IN2[25] | select_2x_4 & IN2[24] | select_n2x_4 & (~ IN2[24]) | select_ne_4 & (~ IN2[25])  );
    wire logic pp_4_26;
    assign pp_4_26 = (select_e_4 & IN2[26] | select_2x_4 & IN2[25] | select_n2x_4 & (~ IN2[25]) | select_ne_4 & (~ IN2[26])  );
    wire logic pp_4_27;
    assign pp_4_27 = (select_e_4 & IN2[27] | select_2x_4 & IN2[26] | select_n2x_4 & (~ IN2[26]) | select_ne_4 & (~ IN2[27])  );
    wire logic pp_4_28;
    assign pp_4_28 = (select_e_4 & IN2[28] | select_2x_4 & IN2[27] | select_n2x_4 & (~ IN2[27]) | select_ne_4 & (~ IN2[28])  );
    wire logic pp_4_29;
    assign pp_4_29 = (select_e_4 & IN2[29] | select_2x_4 & IN2[28] | select_n2x_4 & (~ IN2[28]) | select_ne_4 & (~ IN2[29])  );
    wire logic pp_4_30;
    assign pp_4_30 = (select_e_4 & IN2[30] | select_2x_4 & IN2[29] | select_n2x_4 & (~ IN2[29]) | select_ne_4 & (~ IN2[30])  );
    wire logic pp_4_31;
    assign pp_4_31 = (select_e_4 & IN2[31] | select_2x_4 & IN2[30] | select_n2x_4 & (~ IN2[30]) | select_ne_4 & (~ IN2[31])  );
    wire logic pp_4_32;
    assign pp_4_32 = (select_e_4 & IN2[32] | select_2x_4 & IN2[31] | select_n2x_4 & (~ IN2[31]) | select_ne_4 & (~ IN2[32])  );
    wire logic pp_4_33;
    assign pp_4_33 = (select_e_4 & IN2[33] | select_2x_4 & IN2[32] | select_n2x_4 & (~ IN2[32]) | select_ne_4 & (~ IN2[33])  );
    wire logic pp_4_34;
    assign pp_4_34 = (select_e_4 & IN2[34] | select_2x_4 & IN2[33] | select_n2x_4 & (~ IN2[33]) | select_ne_4 & (~ IN2[34])  );
    wire logic pp_4_35;
    assign pp_4_35 = (select_e_4 & IN2[35] | select_2x_4 & IN2[34] | select_n2x_4 & (~ IN2[34]) | select_ne_4 & (~ IN2[35])  );
    wire logic pp_4_36;
    assign pp_4_36 = (select_e_4 & IN2[36] | select_2x_4 & IN2[35] | select_n2x_4 & (~ IN2[35]) | select_ne_4 & (~ IN2[36])  );
    wire logic pp_4_37;
    assign pp_4_37 = (select_e_4 & IN2[37] | select_2x_4 & IN2[36] | select_n2x_4 & (~ IN2[36]) | select_ne_4 & (~ IN2[37])  );
    wire logic pp_4_38;
    assign pp_4_38 = (select_e_4 & IN2[38] | select_2x_4 & IN2[37] | select_n2x_4 & (~ IN2[37]) | select_ne_4 & (~ IN2[38])  );
    wire logic pp_4_39;
    assign pp_4_39 = (select_e_4 & IN2[39] | select_2x_4 & IN2[38] | select_n2x_4 & (~ IN2[38]) | select_ne_4 & (~ IN2[39])  );
    wire logic pp_4_40;
    assign pp_4_40 = (select_e_4 & IN2[40] | select_2x_4 & IN2[39] | select_n2x_4 & (~ IN2[39]) | select_ne_4 & (~ IN2[40])  );
    wire logic pp_4_41;
    assign pp_4_41 = (select_e_4 & IN2[41] | select_2x_4 & IN2[40] | select_n2x_4 & (~ IN2[40]) | select_ne_4 & (~ IN2[41])  );
    wire logic pp_4_42;
    assign pp_4_42 = (select_e_4 & IN2[42] | select_2x_4 & IN2[41] | select_n2x_4 & (~ IN2[41]) | select_ne_4 & (~ IN2[42])  );
    wire logic pp_4_43;
    assign pp_4_43 = (select_e_4 & IN2[43] | select_2x_4 & IN2[42] | select_n2x_4 & (~ IN2[42]) | select_ne_4 & (~ IN2[43])  );
    wire logic pp_4_44;
    assign pp_4_44 = (select_e_4 & IN2[44] | select_2x_4 & IN2[43] | select_n2x_4 & (~ IN2[43]) | select_ne_4 & (~ IN2[44])  );
    wire logic pp_4_45;
    assign pp_4_45 = (select_e_4 & IN2[45] | select_2x_4 & IN2[44] | select_n2x_4 & (~ IN2[44]) | select_ne_4 & (~ IN2[45])  );
    wire logic pp_4_46;
    assign pp_4_46 = (select_e_4 & IN2[46] | select_2x_4 & IN2[45] | select_n2x_4 & (~ IN2[45]) | select_ne_4 & (~ IN2[46])  );
    wire logic pp_4_47;
    assign pp_4_47 = (select_e_4 & IN2[47] | select_2x_4 & IN2[46] | select_n2x_4 & (~ IN2[46]) | select_ne_4 & (~ IN2[47])  );
    wire logic pp_4_48;
    assign pp_4_48 = (select_e_4 & IN2[48] | select_2x_4 & IN2[47] | select_n2x_4 & (~ IN2[47]) | select_ne_4 & (~ IN2[48])  );
    wire logic pp_4_49;
    assign pp_4_49 = (select_e_4 & IN2[49] | select_2x_4 & IN2[48] | select_n2x_4 & (~ IN2[48]) | select_ne_4 & (~ IN2[49])  );
    wire logic pp_4_50;
    assign pp_4_50 = (select_e_4 & IN2[50] | select_2x_4 & IN2[49] | select_n2x_4 & (~ IN2[49]) | select_ne_4 & (~ IN2[50])  );
    wire logic pp_4_51;
    assign pp_4_51 = (select_e_4 & IN2[51] | select_2x_4 & IN2[50] | select_n2x_4 & (~ IN2[50]) | select_ne_4 & (~ IN2[51])  );
    wire logic pp_4_52;
    assign pp_4_52 = (select_e_4 & IN2[52] | select_2x_4 & IN2[51] | select_n2x_4 & (~ IN2[51]) | select_ne_4 & (~ IN2[52])  );
    wire logic pp_4_53;
    assign pp_4_53 = (select_e_4 & IN2[53] | select_2x_4 & IN2[52] | select_n2x_4 & (~ IN2[52]) | select_ne_4 & (~ IN2[53])  );
    wire logic pp_4_54;
    assign pp_4_54 = (select_e_4 & IN2[54] | select_2x_4 & IN2[53] | select_n2x_4 & (~ IN2[53]) | select_ne_4 & (~ IN2[54])  );
    wire logic pp_4_55;
    assign pp_4_55 = (select_e_4 & IN2[55] | select_2x_4 & IN2[54] | select_n2x_4 & (~ IN2[54]) | select_ne_4 & (~ IN2[55])  );
    wire logic pp_4_56;
    assign pp_4_56 = (select_e_4 & IN2[56] | select_2x_4 & IN2[55] | select_n2x_4 & (~ IN2[55]) | select_ne_4 & (~ IN2[56])  );
    wire logic pp_4_57;
    assign pp_4_57 = (select_e_4 & IN2[57] | select_2x_4 & IN2[56] | select_n2x_4 & (~ IN2[56]) | select_ne_4 & (~ IN2[57])  );
    wire logic pp_4_58;
    assign pp_4_58 = (select_e_4 & IN2[58] | select_2x_4 & IN2[57] | select_n2x_4 & (~ IN2[57]) | select_ne_4 & (~ IN2[58])  );
    wire logic pp_4_59;
    assign pp_4_59 = (select_e_4 & IN2[59] | select_2x_4 & IN2[58] | select_n2x_4 & (~ IN2[58]) | select_ne_4 & (~ IN2[59])  );
    wire logic pp_4_60;
    assign pp_4_60 = (select_e_4 & IN2[60] | select_2x_4 & IN2[59] | select_n2x_4 & (~ IN2[59]) | select_ne_4 & (~ IN2[60])  );
    wire logic pp_4_61;
    assign pp_4_61 = (select_e_4 & IN2[61] | select_2x_4 & IN2[60] | select_n2x_4 & (~ IN2[60]) | select_ne_4 & (~ IN2[61])  );
    wire logic pp_4_62;
    assign pp_4_62 = (select_e_4 & IN2[62] | select_2x_4 & IN2[61] | select_n2x_4 & (~ IN2[61]) | select_ne_4 & (~ IN2[62])  );
    wire logic pp_4_63;
    assign pp_4_63 = (select_e_4 & IN2[63] | select_2x_4 & IN2[62] | select_n2x_4 & (~ IN2[62]) | select_ne_4 & (~ IN2[63])  );
    wire logic pp_4_64;
    assign pp_4_64 = (select_e_4 & IN2[63] | select_2x_4 & IN2[63] | select_n2x_4 & (~ IN2[63]) | select_ne_4 & (~ IN2[63])  );
    wire logic pp_4_65;
    assign pp_4_65 = ~ (select_e_4 & IN2[63] | select_2x_4 & IN2[63] | select_n2x_4 & (~ IN2[63]) | select_ne_4 & (~ IN2[63])  );
    assign tcomp4 = select_ne_4 | select_n2x_4;
    
    // Signed Booth Radix-4 Partial Products Row 6
    wire logic select_e_5, select_ne_5, select_2x_5, tcomp5, select_n2x_5;
    assign select_e_5 = ((~ IN1[11]) & (IN1[10] ^ IN1[9]));
    assign select_ne_5 = IN1[11] &  (IN1[10] ^ IN1[9]);
    assign select_2x_5 = (~ IN1[11]) & IN1[10] & IN1[9];
    assign select_n2x_5 = IN1[11] & (~ IN1[10]) & (~ IN1[9]);
    wire logic pp_5_0;
    assign pp_5_0 = (select_e_5 & IN2[0] | select_2x_5 & 1'b0 | select_n2x_5 & 1'b1 | select_ne_5 & (~ IN2[0])  );
    wire logic pp_5_1;
    assign pp_5_1 = (select_e_5 & IN2[1] | select_2x_5 & IN2[0] | select_n2x_5 & (~ IN2[0]) | select_ne_5 & (~ IN2[1])  );
    wire logic pp_5_2;
    assign pp_5_2 = (select_e_5 & IN2[2] | select_2x_5 & IN2[1] | select_n2x_5 & (~ IN2[1]) | select_ne_5 & (~ IN2[2])  );
    wire logic pp_5_3;
    assign pp_5_3 = (select_e_5 & IN2[3] | select_2x_5 & IN2[2] | select_n2x_5 & (~ IN2[2]) | select_ne_5 & (~ IN2[3])  );
    wire logic pp_5_4;
    assign pp_5_4 = (select_e_5 & IN2[4] | select_2x_5 & IN2[3] | select_n2x_5 & (~ IN2[3]) | select_ne_5 & (~ IN2[4])  );
    wire logic pp_5_5;
    assign pp_5_5 = (select_e_5 & IN2[5] | select_2x_5 & IN2[4] | select_n2x_5 & (~ IN2[4]) | select_ne_5 & (~ IN2[5])  );
    wire logic pp_5_6;
    assign pp_5_6 = (select_e_5 & IN2[6] | select_2x_5 & IN2[5] | select_n2x_5 & (~ IN2[5]) | select_ne_5 & (~ IN2[6])  );
    wire logic pp_5_7;
    assign pp_5_7 = (select_e_5 & IN2[7] | select_2x_5 & IN2[6] | select_n2x_5 & (~ IN2[6]) | select_ne_5 & (~ IN2[7])  );
    wire logic pp_5_8;
    assign pp_5_8 = (select_e_5 & IN2[8] | select_2x_5 & IN2[7] | select_n2x_5 & (~ IN2[7]) | select_ne_5 & (~ IN2[8])  );
    wire logic pp_5_9;
    assign pp_5_9 = (select_e_5 & IN2[9] | select_2x_5 & IN2[8] | select_n2x_5 & (~ IN2[8]) | select_ne_5 & (~ IN2[9])  );
    wire logic pp_5_10;
    assign pp_5_10 = (select_e_5 & IN2[10] | select_2x_5 & IN2[9] | select_n2x_5 & (~ IN2[9]) | select_ne_5 & (~ IN2[10])  );
    wire logic pp_5_11;
    assign pp_5_11 = (select_e_5 & IN2[11] | select_2x_5 & IN2[10] | select_n2x_5 & (~ IN2[10]) | select_ne_5 & (~ IN2[11])  );
    wire logic pp_5_12;
    assign pp_5_12 = (select_e_5 & IN2[12] | select_2x_5 & IN2[11] | select_n2x_5 & (~ IN2[11]) | select_ne_5 & (~ IN2[12])  );
    wire logic pp_5_13;
    assign pp_5_13 = (select_e_5 & IN2[13] | select_2x_5 & IN2[12] | select_n2x_5 & (~ IN2[12]) | select_ne_5 & (~ IN2[13])  );
    wire logic pp_5_14;
    assign pp_5_14 = (select_e_5 & IN2[14] | select_2x_5 & IN2[13] | select_n2x_5 & (~ IN2[13]) | select_ne_5 & (~ IN2[14])  );
    wire logic pp_5_15;
    assign pp_5_15 = (select_e_5 & IN2[15] | select_2x_5 & IN2[14] | select_n2x_5 & (~ IN2[14]) | select_ne_5 & (~ IN2[15])  );
    wire logic pp_5_16;
    assign pp_5_16 = (select_e_5 & IN2[16] | select_2x_5 & IN2[15] | select_n2x_5 & (~ IN2[15]) | select_ne_5 & (~ IN2[16])  );
    wire logic pp_5_17;
    assign pp_5_17 = (select_e_5 & IN2[17] | select_2x_5 & IN2[16] | select_n2x_5 & (~ IN2[16]) | select_ne_5 & (~ IN2[17])  );
    wire logic pp_5_18;
    assign pp_5_18 = (select_e_5 & IN2[18] | select_2x_5 & IN2[17] | select_n2x_5 & (~ IN2[17]) | select_ne_5 & (~ IN2[18])  );
    wire logic pp_5_19;
    assign pp_5_19 = (select_e_5 & IN2[19] | select_2x_5 & IN2[18] | select_n2x_5 & (~ IN2[18]) | select_ne_5 & (~ IN2[19])  );
    wire logic pp_5_20;
    assign pp_5_20 = (select_e_5 & IN2[20] | select_2x_5 & IN2[19] | select_n2x_5 & (~ IN2[19]) | select_ne_5 & (~ IN2[20])  );
    wire logic pp_5_21;
    assign pp_5_21 = (select_e_5 & IN2[21] | select_2x_5 & IN2[20] | select_n2x_5 & (~ IN2[20]) | select_ne_5 & (~ IN2[21])  );
    wire logic pp_5_22;
    assign pp_5_22 = (select_e_5 & IN2[22] | select_2x_5 & IN2[21] | select_n2x_5 & (~ IN2[21]) | select_ne_5 & (~ IN2[22])  );
    wire logic pp_5_23;
    assign pp_5_23 = (select_e_5 & IN2[23] | select_2x_5 & IN2[22] | select_n2x_5 & (~ IN2[22]) | select_ne_5 & (~ IN2[23])  );
    wire logic pp_5_24;
    assign pp_5_24 = (select_e_5 & IN2[24] | select_2x_5 & IN2[23] | select_n2x_5 & (~ IN2[23]) | select_ne_5 & (~ IN2[24])  );
    wire logic pp_5_25;
    assign pp_5_25 = (select_e_5 & IN2[25] | select_2x_5 & IN2[24] | select_n2x_5 & (~ IN2[24]) | select_ne_5 & (~ IN2[25])  );
    wire logic pp_5_26;
    assign pp_5_26 = (select_e_5 & IN2[26] | select_2x_5 & IN2[25] | select_n2x_5 & (~ IN2[25]) | select_ne_5 & (~ IN2[26])  );
    wire logic pp_5_27;
    assign pp_5_27 = (select_e_5 & IN2[27] | select_2x_5 & IN2[26] | select_n2x_5 & (~ IN2[26]) | select_ne_5 & (~ IN2[27])  );
    wire logic pp_5_28;
    assign pp_5_28 = (select_e_5 & IN2[28] | select_2x_5 & IN2[27] | select_n2x_5 & (~ IN2[27]) | select_ne_5 & (~ IN2[28])  );
    wire logic pp_5_29;
    assign pp_5_29 = (select_e_5 & IN2[29] | select_2x_5 & IN2[28] | select_n2x_5 & (~ IN2[28]) | select_ne_5 & (~ IN2[29])  );
    wire logic pp_5_30;
    assign pp_5_30 = (select_e_5 & IN2[30] | select_2x_5 & IN2[29] | select_n2x_5 & (~ IN2[29]) | select_ne_5 & (~ IN2[30])  );
    wire logic pp_5_31;
    assign pp_5_31 = (select_e_5 & IN2[31] | select_2x_5 & IN2[30] | select_n2x_5 & (~ IN2[30]) | select_ne_5 & (~ IN2[31])  );
    wire logic pp_5_32;
    assign pp_5_32 = (select_e_5 & IN2[32] | select_2x_5 & IN2[31] | select_n2x_5 & (~ IN2[31]) | select_ne_5 & (~ IN2[32])  );
    wire logic pp_5_33;
    assign pp_5_33 = (select_e_5 & IN2[33] | select_2x_5 & IN2[32] | select_n2x_5 & (~ IN2[32]) | select_ne_5 & (~ IN2[33])  );
    wire logic pp_5_34;
    assign pp_5_34 = (select_e_5 & IN2[34] | select_2x_5 & IN2[33] | select_n2x_5 & (~ IN2[33]) | select_ne_5 & (~ IN2[34])  );
    wire logic pp_5_35;
    assign pp_5_35 = (select_e_5 & IN2[35] | select_2x_5 & IN2[34] | select_n2x_5 & (~ IN2[34]) | select_ne_5 & (~ IN2[35])  );
    wire logic pp_5_36;
    assign pp_5_36 = (select_e_5 & IN2[36] | select_2x_5 & IN2[35] | select_n2x_5 & (~ IN2[35]) | select_ne_5 & (~ IN2[36])  );
    wire logic pp_5_37;
    assign pp_5_37 = (select_e_5 & IN2[37] | select_2x_5 & IN2[36] | select_n2x_5 & (~ IN2[36]) | select_ne_5 & (~ IN2[37])  );
    wire logic pp_5_38;
    assign pp_5_38 = (select_e_5 & IN2[38] | select_2x_5 & IN2[37] | select_n2x_5 & (~ IN2[37]) | select_ne_5 & (~ IN2[38])  );
    wire logic pp_5_39;
    assign pp_5_39 = (select_e_5 & IN2[39] | select_2x_5 & IN2[38] | select_n2x_5 & (~ IN2[38]) | select_ne_5 & (~ IN2[39])  );
    wire logic pp_5_40;
    assign pp_5_40 = (select_e_5 & IN2[40] | select_2x_5 & IN2[39] | select_n2x_5 & (~ IN2[39]) | select_ne_5 & (~ IN2[40])  );
    wire logic pp_5_41;
    assign pp_5_41 = (select_e_5 & IN2[41] | select_2x_5 & IN2[40] | select_n2x_5 & (~ IN2[40]) | select_ne_5 & (~ IN2[41])  );
    wire logic pp_5_42;
    assign pp_5_42 = (select_e_5 & IN2[42] | select_2x_5 & IN2[41] | select_n2x_5 & (~ IN2[41]) | select_ne_5 & (~ IN2[42])  );
    wire logic pp_5_43;
    assign pp_5_43 = (select_e_5 & IN2[43] | select_2x_5 & IN2[42] | select_n2x_5 & (~ IN2[42]) | select_ne_5 & (~ IN2[43])  );
    wire logic pp_5_44;
    assign pp_5_44 = (select_e_5 & IN2[44] | select_2x_5 & IN2[43] | select_n2x_5 & (~ IN2[43]) | select_ne_5 & (~ IN2[44])  );
    wire logic pp_5_45;
    assign pp_5_45 = (select_e_5 & IN2[45] | select_2x_5 & IN2[44] | select_n2x_5 & (~ IN2[44]) | select_ne_5 & (~ IN2[45])  );
    wire logic pp_5_46;
    assign pp_5_46 = (select_e_5 & IN2[46] | select_2x_5 & IN2[45] | select_n2x_5 & (~ IN2[45]) | select_ne_5 & (~ IN2[46])  );
    wire logic pp_5_47;
    assign pp_5_47 = (select_e_5 & IN2[47] | select_2x_5 & IN2[46] | select_n2x_5 & (~ IN2[46]) | select_ne_5 & (~ IN2[47])  );
    wire logic pp_5_48;
    assign pp_5_48 = (select_e_5 & IN2[48] | select_2x_5 & IN2[47] | select_n2x_5 & (~ IN2[47]) | select_ne_5 & (~ IN2[48])  );
    wire logic pp_5_49;
    assign pp_5_49 = (select_e_5 & IN2[49] | select_2x_5 & IN2[48] | select_n2x_5 & (~ IN2[48]) | select_ne_5 & (~ IN2[49])  );
    wire logic pp_5_50;
    assign pp_5_50 = (select_e_5 & IN2[50] | select_2x_5 & IN2[49] | select_n2x_5 & (~ IN2[49]) | select_ne_5 & (~ IN2[50])  );
    wire logic pp_5_51;
    assign pp_5_51 = (select_e_5 & IN2[51] | select_2x_5 & IN2[50] | select_n2x_5 & (~ IN2[50]) | select_ne_5 & (~ IN2[51])  );
    wire logic pp_5_52;
    assign pp_5_52 = (select_e_5 & IN2[52] | select_2x_5 & IN2[51] | select_n2x_5 & (~ IN2[51]) | select_ne_5 & (~ IN2[52])  );
    wire logic pp_5_53;
    assign pp_5_53 = (select_e_5 & IN2[53] | select_2x_5 & IN2[52] | select_n2x_5 & (~ IN2[52]) | select_ne_5 & (~ IN2[53])  );
    wire logic pp_5_54;
    assign pp_5_54 = (select_e_5 & IN2[54] | select_2x_5 & IN2[53] | select_n2x_5 & (~ IN2[53]) | select_ne_5 & (~ IN2[54])  );
    wire logic pp_5_55;
    assign pp_5_55 = (select_e_5 & IN2[55] | select_2x_5 & IN2[54] | select_n2x_5 & (~ IN2[54]) | select_ne_5 & (~ IN2[55])  );
    wire logic pp_5_56;
    assign pp_5_56 = (select_e_5 & IN2[56] | select_2x_5 & IN2[55] | select_n2x_5 & (~ IN2[55]) | select_ne_5 & (~ IN2[56])  );
    wire logic pp_5_57;
    assign pp_5_57 = (select_e_5 & IN2[57] | select_2x_5 & IN2[56] | select_n2x_5 & (~ IN2[56]) | select_ne_5 & (~ IN2[57])  );
    wire logic pp_5_58;
    assign pp_5_58 = (select_e_5 & IN2[58] | select_2x_5 & IN2[57] | select_n2x_5 & (~ IN2[57]) | select_ne_5 & (~ IN2[58])  );
    wire logic pp_5_59;
    assign pp_5_59 = (select_e_5 & IN2[59] | select_2x_5 & IN2[58] | select_n2x_5 & (~ IN2[58]) | select_ne_5 & (~ IN2[59])  );
    wire logic pp_5_60;
    assign pp_5_60 = (select_e_5 & IN2[60] | select_2x_5 & IN2[59] | select_n2x_5 & (~ IN2[59]) | select_ne_5 & (~ IN2[60])  );
    wire logic pp_5_61;
    assign pp_5_61 = (select_e_5 & IN2[61] | select_2x_5 & IN2[60] | select_n2x_5 & (~ IN2[60]) | select_ne_5 & (~ IN2[61])  );
    wire logic pp_5_62;
    assign pp_5_62 = (select_e_5 & IN2[62] | select_2x_5 & IN2[61] | select_n2x_5 & (~ IN2[61]) | select_ne_5 & (~ IN2[62])  );
    wire logic pp_5_63;
    assign pp_5_63 = (select_e_5 & IN2[63] | select_2x_5 & IN2[62] | select_n2x_5 & (~ IN2[62]) | select_ne_5 & (~ IN2[63])  );
    wire logic pp_5_64;
    assign pp_5_64 = (select_e_5 & IN2[63] | select_2x_5 & IN2[63] | select_n2x_5 & (~ IN2[63]) | select_ne_5 & (~ IN2[63])  );
    wire logic pp_5_65;
    assign pp_5_65 = ~ (select_e_5 & IN2[63] | select_2x_5 & IN2[63] | select_n2x_5 & (~ IN2[63]) | select_ne_5 & (~ IN2[63])  );
    assign tcomp5 = select_ne_5 | select_n2x_5;
    
    // Signed Booth Radix-4 Partial Products Row 7
    wire logic select_e_6, select_ne_6, select_2x_6, tcomp6, select_n2x_6;
    assign select_e_6 = ((~ IN1[13]) & (IN1[12] ^ IN1[11]));
    assign select_ne_6 = IN1[13] &  (IN1[12] ^ IN1[11]);
    assign select_2x_6 = (~ IN1[13]) & IN1[12] & IN1[11];
    assign select_n2x_6 = IN1[13] & (~ IN1[12]) & (~ IN1[11]);
    wire logic pp_6_0;
    assign pp_6_0 = (select_e_6 & IN2[0] | select_2x_6 & 1'b0 | select_n2x_6 & 1'b1 | select_ne_6 & (~ IN2[0])  );
    wire logic pp_6_1;
    assign pp_6_1 = (select_e_6 & IN2[1] | select_2x_6 & IN2[0] | select_n2x_6 & (~ IN2[0]) | select_ne_6 & (~ IN2[1])  );
    wire logic pp_6_2;
    assign pp_6_2 = (select_e_6 & IN2[2] | select_2x_6 & IN2[1] | select_n2x_6 & (~ IN2[1]) | select_ne_6 & (~ IN2[2])  );
    wire logic pp_6_3;
    assign pp_6_3 = (select_e_6 & IN2[3] | select_2x_6 & IN2[2] | select_n2x_6 & (~ IN2[2]) | select_ne_6 & (~ IN2[3])  );
    wire logic pp_6_4;
    assign pp_6_4 = (select_e_6 & IN2[4] | select_2x_6 & IN2[3] | select_n2x_6 & (~ IN2[3]) | select_ne_6 & (~ IN2[4])  );
    wire logic pp_6_5;
    assign pp_6_5 = (select_e_6 & IN2[5] | select_2x_6 & IN2[4] | select_n2x_6 & (~ IN2[4]) | select_ne_6 & (~ IN2[5])  );
    wire logic pp_6_6;
    assign pp_6_6 = (select_e_6 & IN2[6] | select_2x_6 & IN2[5] | select_n2x_6 & (~ IN2[5]) | select_ne_6 & (~ IN2[6])  );
    wire logic pp_6_7;
    assign pp_6_7 = (select_e_6 & IN2[7] | select_2x_6 & IN2[6] | select_n2x_6 & (~ IN2[6]) | select_ne_6 & (~ IN2[7])  );
    wire logic pp_6_8;
    assign pp_6_8 = (select_e_6 & IN2[8] | select_2x_6 & IN2[7] | select_n2x_6 & (~ IN2[7]) | select_ne_6 & (~ IN2[8])  );
    wire logic pp_6_9;
    assign pp_6_9 = (select_e_6 & IN2[9] | select_2x_6 & IN2[8] | select_n2x_6 & (~ IN2[8]) | select_ne_6 & (~ IN2[9])  );
    wire logic pp_6_10;
    assign pp_6_10 = (select_e_6 & IN2[10] | select_2x_6 & IN2[9] | select_n2x_6 & (~ IN2[9]) | select_ne_6 & (~ IN2[10])  );
    wire logic pp_6_11;
    assign pp_6_11 = (select_e_6 & IN2[11] | select_2x_6 & IN2[10] | select_n2x_6 & (~ IN2[10]) | select_ne_6 & (~ IN2[11])  );
    wire logic pp_6_12;
    assign pp_6_12 = (select_e_6 & IN2[12] | select_2x_6 & IN2[11] | select_n2x_6 & (~ IN2[11]) | select_ne_6 & (~ IN2[12])  );
    wire logic pp_6_13;
    assign pp_6_13 = (select_e_6 & IN2[13] | select_2x_6 & IN2[12] | select_n2x_6 & (~ IN2[12]) | select_ne_6 & (~ IN2[13])  );
    wire logic pp_6_14;
    assign pp_6_14 = (select_e_6 & IN2[14] | select_2x_6 & IN2[13] | select_n2x_6 & (~ IN2[13]) | select_ne_6 & (~ IN2[14])  );
    wire logic pp_6_15;
    assign pp_6_15 = (select_e_6 & IN2[15] | select_2x_6 & IN2[14] | select_n2x_6 & (~ IN2[14]) | select_ne_6 & (~ IN2[15])  );
    wire logic pp_6_16;
    assign pp_6_16 = (select_e_6 & IN2[16] | select_2x_6 & IN2[15] | select_n2x_6 & (~ IN2[15]) | select_ne_6 & (~ IN2[16])  );
    wire logic pp_6_17;
    assign pp_6_17 = (select_e_6 & IN2[17] | select_2x_6 & IN2[16] | select_n2x_6 & (~ IN2[16]) | select_ne_6 & (~ IN2[17])  );
    wire logic pp_6_18;
    assign pp_6_18 = (select_e_6 & IN2[18] | select_2x_6 & IN2[17] | select_n2x_6 & (~ IN2[17]) | select_ne_6 & (~ IN2[18])  );
    wire logic pp_6_19;
    assign pp_6_19 = (select_e_6 & IN2[19] | select_2x_6 & IN2[18] | select_n2x_6 & (~ IN2[18]) | select_ne_6 & (~ IN2[19])  );
    wire logic pp_6_20;
    assign pp_6_20 = (select_e_6 & IN2[20] | select_2x_6 & IN2[19] | select_n2x_6 & (~ IN2[19]) | select_ne_6 & (~ IN2[20])  );
    wire logic pp_6_21;
    assign pp_6_21 = (select_e_6 & IN2[21] | select_2x_6 & IN2[20] | select_n2x_6 & (~ IN2[20]) | select_ne_6 & (~ IN2[21])  );
    wire logic pp_6_22;
    assign pp_6_22 = (select_e_6 & IN2[22] | select_2x_6 & IN2[21] | select_n2x_6 & (~ IN2[21]) | select_ne_6 & (~ IN2[22])  );
    wire logic pp_6_23;
    assign pp_6_23 = (select_e_6 & IN2[23] | select_2x_6 & IN2[22] | select_n2x_6 & (~ IN2[22]) | select_ne_6 & (~ IN2[23])  );
    wire logic pp_6_24;
    assign pp_6_24 = (select_e_6 & IN2[24] | select_2x_6 & IN2[23] | select_n2x_6 & (~ IN2[23]) | select_ne_6 & (~ IN2[24])  );
    wire logic pp_6_25;
    assign pp_6_25 = (select_e_6 & IN2[25] | select_2x_6 & IN2[24] | select_n2x_6 & (~ IN2[24]) | select_ne_6 & (~ IN2[25])  );
    wire logic pp_6_26;
    assign pp_6_26 = (select_e_6 & IN2[26] | select_2x_6 & IN2[25] | select_n2x_6 & (~ IN2[25]) | select_ne_6 & (~ IN2[26])  );
    wire logic pp_6_27;
    assign pp_6_27 = (select_e_6 & IN2[27] | select_2x_6 & IN2[26] | select_n2x_6 & (~ IN2[26]) | select_ne_6 & (~ IN2[27])  );
    wire logic pp_6_28;
    assign pp_6_28 = (select_e_6 & IN2[28] | select_2x_6 & IN2[27] | select_n2x_6 & (~ IN2[27]) | select_ne_6 & (~ IN2[28])  );
    wire logic pp_6_29;
    assign pp_6_29 = (select_e_6 & IN2[29] | select_2x_6 & IN2[28] | select_n2x_6 & (~ IN2[28]) | select_ne_6 & (~ IN2[29])  );
    wire logic pp_6_30;
    assign pp_6_30 = (select_e_6 & IN2[30] | select_2x_6 & IN2[29] | select_n2x_6 & (~ IN2[29]) | select_ne_6 & (~ IN2[30])  );
    wire logic pp_6_31;
    assign pp_6_31 = (select_e_6 & IN2[31] | select_2x_6 & IN2[30] | select_n2x_6 & (~ IN2[30]) | select_ne_6 & (~ IN2[31])  );
    wire logic pp_6_32;
    assign pp_6_32 = (select_e_6 & IN2[32] | select_2x_6 & IN2[31] | select_n2x_6 & (~ IN2[31]) | select_ne_6 & (~ IN2[32])  );
    wire logic pp_6_33;
    assign pp_6_33 = (select_e_6 & IN2[33] | select_2x_6 & IN2[32] | select_n2x_6 & (~ IN2[32]) | select_ne_6 & (~ IN2[33])  );
    wire logic pp_6_34;
    assign pp_6_34 = (select_e_6 & IN2[34] | select_2x_6 & IN2[33] | select_n2x_6 & (~ IN2[33]) | select_ne_6 & (~ IN2[34])  );
    wire logic pp_6_35;
    assign pp_6_35 = (select_e_6 & IN2[35] | select_2x_6 & IN2[34] | select_n2x_6 & (~ IN2[34]) | select_ne_6 & (~ IN2[35])  );
    wire logic pp_6_36;
    assign pp_6_36 = (select_e_6 & IN2[36] | select_2x_6 & IN2[35] | select_n2x_6 & (~ IN2[35]) | select_ne_6 & (~ IN2[36])  );
    wire logic pp_6_37;
    assign pp_6_37 = (select_e_6 & IN2[37] | select_2x_6 & IN2[36] | select_n2x_6 & (~ IN2[36]) | select_ne_6 & (~ IN2[37])  );
    wire logic pp_6_38;
    assign pp_6_38 = (select_e_6 & IN2[38] | select_2x_6 & IN2[37] | select_n2x_6 & (~ IN2[37]) | select_ne_6 & (~ IN2[38])  );
    wire logic pp_6_39;
    assign pp_6_39 = (select_e_6 & IN2[39] | select_2x_6 & IN2[38] | select_n2x_6 & (~ IN2[38]) | select_ne_6 & (~ IN2[39])  );
    wire logic pp_6_40;
    assign pp_6_40 = (select_e_6 & IN2[40] | select_2x_6 & IN2[39] | select_n2x_6 & (~ IN2[39]) | select_ne_6 & (~ IN2[40])  );
    wire logic pp_6_41;
    assign pp_6_41 = (select_e_6 & IN2[41] | select_2x_6 & IN2[40] | select_n2x_6 & (~ IN2[40]) | select_ne_6 & (~ IN2[41])  );
    wire logic pp_6_42;
    assign pp_6_42 = (select_e_6 & IN2[42] | select_2x_6 & IN2[41] | select_n2x_6 & (~ IN2[41]) | select_ne_6 & (~ IN2[42])  );
    wire logic pp_6_43;
    assign pp_6_43 = (select_e_6 & IN2[43] | select_2x_6 & IN2[42] | select_n2x_6 & (~ IN2[42]) | select_ne_6 & (~ IN2[43])  );
    wire logic pp_6_44;
    assign pp_6_44 = (select_e_6 & IN2[44] | select_2x_6 & IN2[43] | select_n2x_6 & (~ IN2[43]) | select_ne_6 & (~ IN2[44])  );
    wire logic pp_6_45;
    assign pp_6_45 = (select_e_6 & IN2[45] | select_2x_6 & IN2[44] | select_n2x_6 & (~ IN2[44]) | select_ne_6 & (~ IN2[45])  );
    wire logic pp_6_46;
    assign pp_6_46 = (select_e_6 & IN2[46] | select_2x_6 & IN2[45] | select_n2x_6 & (~ IN2[45]) | select_ne_6 & (~ IN2[46])  );
    wire logic pp_6_47;
    assign pp_6_47 = (select_e_6 & IN2[47] | select_2x_6 & IN2[46] | select_n2x_6 & (~ IN2[46]) | select_ne_6 & (~ IN2[47])  );
    wire logic pp_6_48;
    assign pp_6_48 = (select_e_6 & IN2[48] | select_2x_6 & IN2[47] | select_n2x_6 & (~ IN2[47]) | select_ne_6 & (~ IN2[48])  );
    wire logic pp_6_49;
    assign pp_6_49 = (select_e_6 & IN2[49] | select_2x_6 & IN2[48] | select_n2x_6 & (~ IN2[48]) | select_ne_6 & (~ IN2[49])  );
    wire logic pp_6_50;
    assign pp_6_50 = (select_e_6 & IN2[50] | select_2x_6 & IN2[49] | select_n2x_6 & (~ IN2[49]) | select_ne_6 & (~ IN2[50])  );
    wire logic pp_6_51;
    assign pp_6_51 = (select_e_6 & IN2[51] | select_2x_6 & IN2[50] | select_n2x_6 & (~ IN2[50]) | select_ne_6 & (~ IN2[51])  );
    wire logic pp_6_52;
    assign pp_6_52 = (select_e_6 & IN2[52] | select_2x_6 & IN2[51] | select_n2x_6 & (~ IN2[51]) | select_ne_6 & (~ IN2[52])  );
    wire logic pp_6_53;
    assign pp_6_53 = (select_e_6 & IN2[53] | select_2x_6 & IN2[52] | select_n2x_6 & (~ IN2[52]) | select_ne_6 & (~ IN2[53])  );
    wire logic pp_6_54;
    assign pp_6_54 = (select_e_6 & IN2[54] | select_2x_6 & IN2[53] | select_n2x_6 & (~ IN2[53]) | select_ne_6 & (~ IN2[54])  );
    wire logic pp_6_55;
    assign pp_6_55 = (select_e_6 & IN2[55] | select_2x_6 & IN2[54] | select_n2x_6 & (~ IN2[54]) | select_ne_6 & (~ IN2[55])  );
    wire logic pp_6_56;
    assign pp_6_56 = (select_e_6 & IN2[56] | select_2x_6 & IN2[55] | select_n2x_6 & (~ IN2[55]) | select_ne_6 & (~ IN2[56])  );
    wire logic pp_6_57;
    assign pp_6_57 = (select_e_6 & IN2[57] | select_2x_6 & IN2[56] | select_n2x_6 & (~ IN2[56]) | select_ne_6 & (~ IN2[57])  );
    wire logic pp_6_58;
    assign pp_6_58 = (select_e_6 & IN2[58] | select_2x_6 & IN2[57] | select_n2x_6 & (~ IN2[57]) | select_ne_6 & (~ IN2[58])  );
    wire logic pp_6_59;
    assign pp_6_59 = (select_e_6 & IN2[59] | select_2x_6 & IN2[58] | select_n2x_6 & (~ IN2[58]) | select_ne_6 & (~ IN2[59])  );
    wire logic pp_6_60;
    assign pp_6_60 = (select_e_6 & IN2[60] | select_2x_6 & IN2[59] | select_n2x_6 & (~ IN2[59]) | select_ne_6 & (~ IN2[60])  );
    wire logic pp_6_61;
    assign pp_6_61 = (select_e_6 & IN2[61] | select_2x_6 & IN2[60] | select_n2x_6 & (~ IN2[60]) | select_ne_6 & (~ IN2[61])  );
    wire logic pp_6_62;
    assign pp_6_62 = (select_e_6 & IN2[62] | select_2x_6 & IN2[61] | select_n2x_6 & (~ IN2[61]) | select_ne_6 & (~ IN2[62])  );
    wire logic pp_6_63;
    assign pp_6_63 = (select_e_6 & IN2[63] | select_2x_6 & IN2[62] | select_n2x_6 & (~ IN2[62]) | select_ne_6 & (~ IN2[63])  );
    wire logic pp_6_64;
    assign pp_6_64 = (select_e_6 & IN2[63] | select_2x_6 & IN2[63] | select_n2x_6 & (~ IN2[63]) | select_ne_6 & (~ IN2[63])  );
    wire logic pp_6_65;
    assign pp_6_65 = ~ (select_e_6 & IN2[63] | select_2x_6 & IN2[63] | select_n2x_6 & (~ IN2[63]) | select_ne_6 & (~ IN2[63])  );
    assign tcomp6 = select_ne_6 | select_n2x_6;
    
    // Signed Booth Radix-4 Partial Products Row 8
    wire logic select_e_7, select_ne_7, select_2x_7, tcomp7, select_n2x_7;
    assign select_e_7 = ((~ IN1[15]) & (IN1[14] ^ IN1[13]));
    assign select_ne_7 = IN1[15] &  (IN1[14] ^ IN1[13]);
    assign select_2x_7 = (~ IN1[15]) & IN1[14] & IN1[13];
    assign select_n2x_7 = IN1[15] & (~ IN1[14]) & (~ IN1[13]);
    wire logic pp_7_0;
    assign pp_7_0 = (select_e_7 & IN2[0] | select_2x_7 & 1'b0 | select_n2x_7 & 1'b1 | select_ne_7 & (~ IN2[0])  );
    wire logic pp_7_1;
    assign pp_7_1 = (select_e_7 & IN2[1] | select_2x_7 & IN2[0] | select_n2x_7 & (~ IN2[0]) | select_ne_7 & (~ IN2[1])  );
    wire logic pp_7_2;
    assign pp_7_2 = (select_e_7 & IN2[2] | select_2x_7 & IN2[1] | select_n2x_7 & (~ IN2[1]) | select_ne_7 & (~ IN2[2])  );
    wire logic pp_7_3;
    assign pp_7_3 = (select_e_7 & IN2[3] | select_2x_7 & IN2[2] | select_n2x_7 & (~ IN2[2]) | select_ne_7 & (~ IN2[3])  );
    wire logic pp_7_4;
    assign pp_7_4 = (select_e_7 & IN2[4] | select_2x_7 & IN2[3] | select_n2x_7 & (~ IN2[3]) | select_ne_7 & (~ IN2[4])  );
    wire logic pp_7_5;
    assign pp_7_5 = (select_e_7 & IN2[5] | select_2x_7 & IN2[4] | select_n2x_7 & (~ IN2[4]) | select_ne_7 & (~ IN2[5])  );
    wire logic pp_7_6;
    assign pp_7_6 = (select_e_7 & IN2[6] | select_2x_7 & IN2[5] | select_n2x_7 & (~ IN2[5]) | select_ne_7 & (~ IN2[6])  );
    wire logic pp_7_7;
    assign pp_7_7 = (select_e_7 & IN2[7] | select_2x_7 & IN2[6] | select_n2x_7 & (~ IN2[6]) | select_ne_7 & (~ IN2[7])  );
    wire logic pp_7_8;
    assign pp_7_8 = (select_e_7 & IN2[8] | select_2x_7 & IN2[7] | select_n2x_7 & (~ IN2[7]) | select_ne_7 & (~ IN2[8])  );
    wire logic pp_7_9;
    assign pp_7_9 = (select_e_7 & IN2[9] | select_2x_7 & IN2[8] | select_n2x_7 & (~ IN2[8]) | select_ne_7 & (~ IN2[9])  );
    wire logic pp_7_10;
    assign pp_7_10 = (select_e_7 & IN2[10] | select_2x_7 & IN2[9] | select_n2x_7 & (~ IN2[9]) | select_ne_7 & (~ IN2[10])  );
    wire logic pp_7_11;
    assign pp_7_11 = (select_e_7 & IN2[11] | select_2x_7 & IN2[10] | select_n2x_7 & (~ IN2[10]) | select_ne_7 & (~ IN2[11])  );
    wire logic pp_7_12;
    assign pp_7_12 = (select_e_7 & IN2[12] | select_2x_7 & IN2[11] | select_n2x_7 & (~ IN2[11]) | select_ne_7 & (~ IN2[12])  );
    wire logic pp_7_13;
    assign pp_7_13 = (select_e_7 & IN2[13] | select_2x_7 & IN2[12] | select_n2x_7 & (~ IN2[12]) | select_ne_7 & (~ IN2[13])  );
    wire logic pp_7_14;
    assign pp_7_14 = (select_e_7 & IN2[14] | select_2x_7 & IN2[13] | select_n2x_7 & (~ IN2[13]) | select_ne_7 & (~ IN2[14])  );
    wire logic pp_7_15;
    assign pp_7_15 = (select_e_7 & IN2[15] | select_2x_7 & IN2[14] | select_n2x_7 & (~ IN2[14]) | select_ne_7 & (~ IN2[15])  );
    wire logic pp_7_16;
    assign pp_7_16 = (select_e_7 & IN2[16] | select_2x_7 & IN2[15] | select_n2x_7 & (~ IN2[15]) | select_ne_7 & (~ IN2[16])  );
    wire logic pp_7_17;
    assign pp_7_17 = (select_e_7 & IN2[17] | select_2x_7 & IN2[16] | select_n2x_7 & (~ IN2[16]) | select_ne_7 & (~ IN2[17])  );
    wire logic pp_7_18;
    assign pp_7_18 = (select_e_7 & IN2[18] | select_2x_7 & IN2[17] | select_n2x_7 & (~ IN2[17]) | select_ne_7 & (~ IN2[18])  );
    wire logic pp_7_19;
    assign pp_7_19 = (select_e_7 & IN2[19] | select_2x_7 & IN2[18] | select_n2x_7 & (~ IN2[18]) | select_ne_7 & (~ IN2[19])  );
    wire logic pp_7_20;
    assign pp_7_20 = (select_e_7 & IN2[20] | select_2x_7 & IN2[19] | select_n2x_7 & (~ IN2[19]) | select_ne_7 & (~ IN2[20])  );
    wire logic pp_7_21;
    assign pp_7_21 = (select_e_7 & IN2[21] | select_2x_7 & IN2[20] | select_n2x_7 & (~ IN2[20]) | select_ne_7 & (~ IN2[21])  );
    wire logic pp_7_22;
    assign pp_7_22 = (select_e_7 & IN2[22] | select_2x_7 & IN2[21] | select_n2x_7 & (~ IN2[21]) | select_ne_7 & (~ IN2[22])  );
    wire logic pp_7_23;
    assign pp_7_23 = (select_e_7 & IN2[23] | select_2x_7 & IN2[22] | select_n2x_7 & (~ IN2[22]) | select_ne_7 & (~ IN2[23])  );
    wire logic pp_7_24;
    assign pp_7_24 = (select_e_7 & IN2[24] | select_2x_7 & IN2[23] | select_n2x_7 & (~ IN2[23]) | select_ne_7 & (~ IN2[24])  );
    wire logic pp_7_25;
    assign pp_7_25 = (select_e_7 & IN2[25] | select_2x_7 & IN2[24] | select_n2x_7 & (~ IN2[24]) | select_ne_7 & (~ IN2[25])  );
    wire logic pp_7_26;
    assign pp_7_26 = (select_e_7 & IN2[26] | select_2x_7 & IN2[25] | select_n2x_7 & (~ IN2[25]) | select_ne_7 & (~ IN2[26])  );
    wire logic pp_7_27;
    assign pp_7_27 = (select_e_7 & IN2[27] | select_2x_7 & IN2[26] | select_n2x_7 & (~ IN2[26]) | select_ne_7 & (~ IN2[27])  );
    wire logic pp_7_28;
    assign pp_7_28 = (select_e_7 & IN2[28] | select_2x_7 & IN2[27] | select_n2x_7 & (~ IN2[27]) | select_ne_7 & (~ IN2[28])  );
    wire logic pp_7_29;
    assign pp_7_29 = (select_e_7 & IN2[29] | select_2x_7 & IN2[28] | select_n2x_7 & (~ IN2[28]) | select_ne_7 & (~ IN2[29])  );
    wire logic pp_7_30;
    assign pp_7_30 = (select_e_7 & IN2[30] | select_2x_7 & IN2[29] | select_n2x_7 & (~ IN2[29]) | select_ne_7 & (~ IN2[30])  );
    wire logic pp_7_31;
    assign pp_7_31 = (select_e_7 & IN2[31] | select_2x_7 & IN2[30] | select_n2x_7 & (~ IN2[30]) | select_ne_7 & (~ IN2[31])  );
    wire logic pp_7_32;
    assign pp_7_32 = (select_e_7 & IN2[32] | select_2x_7 & IN2[31] | select_n2x_7 & (~ IN2[31]) | select_ne_7 & (~ IN2[32])  );
    wire logic pp_7_33;
    assign pp_7_33 = (select_e_7 & IN2[33] | select_2x_7 & IN2[32] | select_n2x_7 & (~ IN2[32]) | select_ne_7 & (~ IN2[33])  );
    wire logic pp_7_34;
    assign pp_7_34 = (select_e_7 & IN2[34] | select_2x_7 & IN2[33] | select_n2x_7 & (~ IN2[33]) | select_ne_7 & (~ IN2[34])  );
    wire logic pp_7_35;
    assign pp_7_35 = (select_e_7 & IN2[35] | select_2x_7 & IN2[34] | select_n2x_7 & (~ IN2[34]) | select_ne_7 & (~ IN2[35])  );
    wire logic pp_7_36;
    assign pp_7_36 = (select_e_7 & IN2[36] | select_2x_7 & IN2[35] | select_n2x_7 & (~ IN2[35]) | select_ne_7 & (~ IN2[36])  );
    wire logic pp_7_37;
    assign pp_7_37 = (select_e_7 & IN2[37] | select_2x_7 & IN2[36] | select_n2x_7 & (~ IN2[36]) | select_ne_7 & (~ IN2[37])  );
    wire logic pp_7_38;
    assign pp_7_38 = (select_e_7 & IN2[38] | select_2x_7 & IN2[37] | select_n2x_7 & (~ IN2[37]) | select_ne_7 & (~ IN2[38])  );
    wire logic pp_7_39;
    assign pp_7_39 = (select_e_7 & IN2[39] | select_2x_7 & IN2[38] | select_n2x_7 & (~ IN2[38]) | select_ne_7 & (~ IN2[39])  );
    wire logic pp_7_40;
    assign pp_7_40 = (select_e_7 & IN2[40] | select_2x_7 & IN2[39] | select_n2x_7 & (~ IN2[39]) | select_ne_7 & (~ IN2[40])  );
    wire logic pp_7_41;
    assign pp_7_41 = (select_e_7 & IN2[41] | select_2x_7 & IN2[40] | select_n2x_7 & (~ IN2[40]) | select_ne_7 & (~ IN2[41])  );
    wire logic pp_7_42;
    assign pp_7_42 = (select_e_7 & IN2[42] | select_2x_7 & IN2[41] | select_n2x_7 & (~ IN2[41]) | select_ne_7 & (~ IN2[42])  );
    wire logic pp_7_43;
    assign pp_7_43 = (select_e_7 & IN2[43] | select_2x_7 & IN2[42] | select_n2x_7 & (~ IN2[42]) | select_ne_7 & (~ IN2[43])  );
    wire logic pp_7_44;
    assign pp_7_44 = (select_e_7 & IN2[44] | select_2x_7 & IN2[43] | select_n2x_7 & (~ IN2[43]) | select_ne_7 & (~ IN2[44])  );
    wire logic pp_7_45;
    assign pp_7_45 = (select_e_7 & IN2[45] | select_2x_7 & IN2[44] | select_n2x_7 & (~ IN2[44]) | select_ne_7 & (~ IN2[45])  );
    wire logic pp_7_46;
    assign pp_7_46 = (select_e_7 & IN2[46] | select_2x_7 & IN2[45] | select_n2x_7 & (~ IN2[45]) | select_ne_7 & (~ IN2[46])  );
    wire logic pp_7_47;
    assign pp_7_47 = (select_e_7 & IN2[47] | select_2x_7 & IN2[46] | select_n2x_7 & (~ IN2[46]) | select_ne_7 & (~ IN2[47])  );
    wire logic pp_7_48;
    assign pp_7_48 = (select_e_7 & IN2[48] | select_2x_7 & IN2[47] | select_n2x_7 & (~ IN2[47]) | select_ne_7 & (~ IN2[48])  );
    wire logic pp_7_49;
    assign pp_7_49 = (select_e_7 & IN2[49] | select_2x_7 & IN2[48] | select_n2x_7 & (~ IN2[48]) | select_ne_7 & (~ IN2[49])  );
    wire logic pp_7_50;
    assign pp_7_50 = (select_e_7 & IN2[50] | select_2x_7 & IN2[49] | select_n2x_7 & (~ IN2[49]) | select_ne_7 & (~ IN2[50])  );
    wire logic pp_7_51;
    assign pp_7_51 = (select_e_7 & IN2[51] | select_2x_7 & IN2[50] | select_n2x_7 & (~ IN2[50]) | select_ne_7 & (~ IN2[51])  );
    wire logic pp_7_52;
    assign pp_7_52 = (select_e_7 & IN2[52] | select_2x_7 & IN2[51] | select_n2x_7 & (~ IN2[51]) | select_ne_7 & (~ IN2[52])  );
    wire logic pp_7_53;
    assign pp_7_53 = (select_e_7 & IN2[53] | select_2x_7 & IN2[52] | select_n2x_7 & (~ IN2[52]) | select_ne_7 & (~ IN2[53])  );
    wire logic pp_7_54;
    assign pp_7_54 = (select_e_7 & IN2[54] | select_2x_7 & IN2[53] | select_n2x_7 & (~ IN2[53]) | select_ne_7 & (~ IN2[54])  );
    wire logic pp_7_55;
    assign pp_7_55 = (select_e_7 & IN2[55] | select_2x_7 & IN2[54] | select_n2x_7 & (~ IN2[54]) | select_ne_7 & (~ IN2[55])  );
    wire logic pp_7_56;
    assign pp_7_56 = (select_e_7 & IN2[56] | select_2x_7 & IN2[55] | select_n2x_7 & (~ IN2[55]) | select_ne_7 & (~ IN2[56])  );
    wire logic pp_7_57;
    assign pp_7_57 = (select_e_7 & IN2[57] | select_2x_7 & IN2[56] | select_n2x_7 & (~ IN2[56]) | select_ne_7 & (~ IN2[57])  );
    wire logic pp_7_58;
    assign pp_7_58 = (select_e_7 & IN2[58] | select_2x_7 & IN2[57] | select_n2x_7 & (~ IN2[57]) | select_ne_7 & (~ IN2[58])  );
    wire logic pp_7_59;
    assign pp_7_59 = (select_e_7 & IN2[59] | select_2x_7 & IN2[58] | select_n2x_7 & (~ IN2[58]) | select_ne_7 & (~ IN2[59])  );
    wire logic pp_7_60;
    assign pp_7_60 = (select_e_7 & IN2[60] | select_2x_7 & IN2[59] | select_n2x_7 & (~ IN2[59]) | select_ne_7 & (~ IN2[60])  );
    wire logic pp_7_61;
    assign pp_7_61 = (select_e_7 & IN2[61] | select_2x_7 & IN2[60] | select_n2x_7 & (~ IN2[60]) | select_ne_7 & (~ IN2[61])  );
    wire logic pp_7_62;
    assign pp_7_62 = (select_e_7 & IN2[62] | select_2x_7 & IN2[61] | select_n2x_7 & (~ IN2[61]) | select_ne_7 & (~ IN2[62])  );
    wire logic pp_7_63;
    assign pp_7_63 = (select_e_7 & IN2[63] | select_2x_7 & IN2[62] | select_n2x_7 & (~ IN2[62]) | select_ne_7 & (~ IN2[63])  );
    wire logic pp_7_64;
    assign pp_7_64 = (select_e_7 & IN2[63] | select_2x_7 & IN2[63] | select_n2x_7 & (~ IN2[63]) | select_ne_7 & (~ IN2[63])  );
    wire logic pp_7_65;
    assign pp_7_65 = ~ (select_e_7 & IN2[63] | select_2x_7 & IN2[63] | select_n2x_7 & (~ IN2[63]) | select_ne_7 & (~ IN2[63])  );
    assign tcomp7 = select_ne_7 | select_n2x_7;
    
    // Signed Booth Radix-4 Partial Products Row 9
    wire logic select_e_8, select_ne_8, select_2x_8, tcomp8, select_n2x_8;
    assign select_e_8 = ((~ IN1[17]) & (IN1[16] ^ IN1[15]));
    assign select_ne_8 = IN1[17] &  (IN1[16] ^ IN1[15]);
    assign select_2x_8 = (~ IN1[17]) & IN1[16] & IN1[15];
    assign select_n2x_8 = IN1[17] & (~ IN1[16]) & (~ IN1[15]);
    wire logic pp_8_0;
    assign pp_8_0 = (select_e_8 & IN2[0] | select_2x_8 & 1'b0 | select_n2x_8 & 1'b1 | select_ne_8 & (~ IN2[0])  );
    wire logic pp_8_1;
    assign pp_8_1 = (select_e_8 & IN2[1] | select_2x_8 & IN2[0] | select_n2x_8 & (~ IN2[0]) | select_ne_8 & (~ IN2[1])  );
    wire logic pp_8_2;
    assign pp_8_2 = (select_e_8 & IN2[2] | select_2x_8 & IN2[1] | select_n2x_8 & (~ IN2[1]) | select_ne_8 & (~ IN2[2])  );
    wire logic pp_8_3;
    assign pp_8_3 = (select_e_8 & IN2[3] | select_2x_8 & IN2[2] | select_n2x_8 & (~ IN2[2]) | select_ne_8 & (~ IN2[3])  );
    wire logic pp_8_4;
    assign pp_8_4 = (select_e_8 & IN2[4] | select_2x_8 & IN2[3] | select_n2x_8 & (~ IN2[3]) | select_ne_8 & (~ IN2[4])  );
    wire logic pp_8_5;
    assign pp_8_5 = (select_e_8 & IN2[5] | select_2x_8 & IN2[4] | select_n2x_8 & (~ IN2[4]) | select_ne_8 & (~ IN2[5])  );
    wire logic pp_8_6;
    assign pp_8_6 = (select_e_8 & IN2[6] | select_2x_8 & IN2[5] | select_n2x_8 & (~ IN2[5]) | select_ne_8 & (~ IN2[6])  );
    wire logic pp_8_7;
    assign pp_8_7 = (select_e_8 & IN2[7] | select_2x_8 & IN2[6] | select_n2x_8 & (~ IN2[6]) | select_ne_8 & (~ IN2[7])  );
    wire logic pp_8_8;
    assign pp_8_8 = (select_e_8 & IN2[8] | select_2x_8 & IN2[7] | select_n2x_8 & (~ IN2[7]) | select_ne_8 & (~ IN2[8])  );
    wire logic pp_8_9;
    assign pp_8_9 = (select_e_8 & IN2[9] | select_2x_8 & IN2[8] | select_n2x_8 & (~ IN2[8]) | select_ne_8 & (~ IN2[9])  );
    wire logic pp_8_10;
    assign pp_8_10 = (select_e_8 & IN2[10] | select_2x_8 & IN2[9] | select_n2x_8 & (~ IN2[9]) | select_ne_8 & (~ IN2[10])  );
    wire logic pp_8_11;
    assign pp_8_11 = (select_e_8 & IN2[11] | select_2x_8 & IN2[10] | select_n2x_8 & (~ IN2[10]) | select_ne_8 & (~ IN2[11])  );
    wire logic pp_8_12;
    assign pp_8_12 = (select_e_8 & IN2[12] | select_2x_8 & IN2[11] | select_n2x_8 & (~ IN2[11]) | select_ne_8 & (~ IN2[12])  );
    wire logic pp_8_13;
    assign pp_8_13 = (select_e_8 & IN2[13] | select_2x_8 & IN2[12] | select_n2x_8 & (~ IN2[12]) | select_ne_8 & (~ IN2[13])  );
    wire logic pp_8_14;
    assign pp_8_14 = (select_e_8 & IN2[14] | select_2x_8 & IN2[13] | select_n2x_8 & (~ IN2[13]) | select_ne_8 & (~ IN2[14])  );
    wire logic pp_8_15;
    assign pp_8_15 = (select_e_8 & IN2[15] | select_2x_8 & IN2[14] | select_n2x_8 & (~ IN2[14]) | select_ne_8 & (~ IN2[15])  );
    wire logic pp_8_16;
    assign pp_8_16 = (select_e_8 & IN2[16] | select_2x_8 & IN2[15] | select_n2x_8 & (~ IN2[15]) | select_ne_8 & (~ IN2[16])  );
    wire logic pp_8_17;
    assign pp_8_17 = (select_e_8 & IN2[17] | select_2x_8 & IN2[16] | select_n2x_8 & (~ IN2[16]) | select_ne_8 & (~ IN2[17])  );
    wire logic pp_8_18;
    assign pp_8_18 = (select_e_8 & IN2[18] | select_2x_8 & IN2[17] | select_n2x_8 & (~ IN2[17]) | select_ne_8 & (~ IN2[18])  );
    wire logic pp_8_19;
    assign pp_8_19 = (select_e_8 & IN2[19] | select_2x_8 & IN2[18] | select_n2x_8 & (~ IN2[18]) | select_ne_8 & (~ IN2[19])  );
    wire logic pp_8_20;
    assign pp_8_20 = (select_e_8 & IN2[20] | select_2x_8 & IN2[19] | select_n2x_8 & (~ IN2[19]) | select_ne_8 & (~ IN2[20])  );
    wire logic pp_8_21;
    assign pp_8_21 = (select_e_8 & IN2[21] | select_2x_8 & IN2[20] | select_n2x_8 & (~ IN2[20]) | select_ne_8 & (~ IN2[21])  );
    wire logic pp_8_22;
    assign pp_8_22 = (select_e_8 & IN2[22] | select_2x_8 & IN2[21] | select_n2x_8 & (~ IN2[21]) | select_ne_8 & (~ IN2[22])  );
    wire logic pp_8_23;
    assign pp_8_23 = (select_e_8 & IN2[23] | select_2x_8 & IN2[22] | select_n2x_8 & (~ IN2[22]) | select_ne_8 & (~ IN2[23])  );
    wire logic pp_8_24;
    assign pp_8_24 = (select_e_8 & IN2[24] | select_2x_8 & IN2[23] | select_n2x_8 & (~ IN2[23]) | select_ne_8 & (~ IN2[24])  );
    wire logic pp_8_25;
    assign pp_8_25 = (select_e_8 & IN2[25] | select_2x_8 & IN2[24] | select_n2x_8 & (~ IN2[24]) | select_ne_8 & (~ IN2[25])  );
    wire logic pp_8_26;
    assign pp_8_26 = (select_e_8 & IN2[26] | select_2x_8 & IN2[25] | select_n2x_8 & (~ IN2[25]) | select_ne_8 & (~ IN2[26])  );
    wire logic pp_8_27;
    assign pp_8_27 = (select_e_8 & IN2[27] | select_2x_8 & IN2[26] | select_n2x_8 & (~ IN2[26]) | select_ne_8 & (~ IN2[27])  );
    wire logic pp_8_28;
    assign pp_8_28 = (select_e_8 & IN2[28] | select_2x_8 & IN2[27] | select_n2x_8 & (~ IN2[27]) | select_ne_8 & (~ IN2[28])  );
    wire logic pp_8_29;
    assign pp_8_29 = (select_e_8 & IN2[29] | select_2x_8 & IN2[28] | select_n2x_8 & (~ IN2[28]) | select_ne_8 & (~ IN2[29])  );
    wire logic pp_8_30;
    assign pp_8_30 = (select_e_8 & IN2[30] | select_2x_8 & IN2[29] | select_n2x_8 & (~ IN2[29]) | select_ne_8 & (~ IN2[30])  );
    wire logic pp_8_31;
    assign pp_8_31 = (select_e_8 & IN2[31] | select_2x_8 & IN2[30] | select_n2x_8 & (~ IN2[30]) | select_ne_8 & (~ IN2[31])  );
    wire logic pp_8_32;
    assign pp_8_32 = (select_e_8 & IN2[32] | select_2x_8 & IN2[31] | select_n2x_8 & (~ IN2[31]) | select_ne_8 & (~ IN2[32])  );
    wire logic pp_8_33;
    assign pp_8_33 = (select_e_8 & IN2[33] | select_2x_8 & IN2[32] | select_n2x_8 & (~ IN2[32]) | select_ne_8 & (~ IN2[33])  );
    wire logic pp_8_34;
    assign pp_8_34 = (select_e_8 & IN2[34] | select_2x_8 & IN2[33] | select_n2x_8 & (~ IN2[33]) | select_ne_8 & (~ IN2[34])  );
    wire logic pp_8_35;
    assign pp_8_35 = (select_e_8 & IN2[35] | select_2x_8 & IN2[34] | select_n2x_8 & (~ IN2[34]) | select_ne_8 & (~ IN2[35])  );
    wire logic pp_8_36;
    assign pp_8_36 = (select_e_8 & IN2[36] | select_2x_8 & IN2[35] | select_n2x_8 & (~ IN2[35]) | select_ne_8 & (~ IN2[36])  );
    wire logic pp_8_37;
    assign pp_8_37 = (select_e_8 & IN2[37] | select_2x_8 & IN2[36] | select_n2x_8 & (~ IN2[36]) | select_ne_8 & (~ IN2[37])  );
    wire logic pp_8_38;
    assign pp_8_38 = (select_e_8 & IN2[38] | select_2x_8 & IN2[37] | select_n2x_8 & (~ IN2[37]) | select_ne_8 & (~ IN2[38])  );
    wire logic pp_8_39;
    assign pp_8_39 = (select_e_8 & IN2[39] | select_2x_8 & IN2[38] | select_n2x_8 & (~ IN2[38]) | select_ne_8 & (~ IN2[39])  );
    wire logic pp_8_40;
    assign pp_8_40 = (select_e_8 & IN2[40] | select_2x_8 & IN2[39] | select_n2x_8 & (~ IN2[39]) | select_ne_8 & (~ IN2[40])  );
    wire logic pp_8_41;
    assign pp_8_41 = (select_e_8 & IN2[41] | select_2x_8 & IN2[40] | select_n2x_8 & (~ IN2[40]) | select_ne_8 & (~ IN2[41])  );
    wire logic pp_8_42;
    assign pp_8_42 = (select_e_8 & IN2[42] | select_2x_8 & IN2[41] | select_n2x_8 & (~ IN2[41]) | select_ne_8 & (~ IN2[42])  );
    wire logic pp_8_43;
    assign pp_8_43 = (select_e_8 & IN2[43] | select_2x_8 & IN2[42] | select_n2x_8 & (~ IN2[42]) | select_ne_8 & (~ IN2[43])  );
    wire logic pp_8_44;
    assign pp_8_44 = (select_e_8 & IN2[44] | select_2x_8 & IN2[43] | select_n2x_8 & (~ IN2[43]) | select_ne_8 & (~ IN2[44])  );
    wire logic pp_8_45;
    assign pp_8_45 = (select_e_8 & IN2[45] | select_2x_8 & IN2[44] | select_n2x_8 & (~ IN2[44]) | select_ne_8 & (~ IN2[45])  );
    wire logic pp_8_46;
    assign pp_8_46 = (select_e_8 & IN2[46] | select_2x_8 & IN2[45] | select_n2x_8 & (~ IN2[45]) | select_ne_8 & (~ IN2[46])  );
    wire logic pp_8_47;
    assign pp_8_47 = (select_e_8 & IN2[47] | select_2x_8 & IN2[46] | select_n2x_8 & (~ IN2[46]) | select_ne_8 & (~ IN2[47])  );
    wire logic pp_8_48;
    assign pp_8_48 = (select_e_8 & IN2[48] | select_2x_8 & IN2[47] | select_n2x_8 & (~ IN2[47]) | select_ne_8 & (~ IN2[48])  );
    wire logic pp_8_49;
    assign pp_8_49 = (select_e_8 & IN2[49] | select_2x_8 & IN2[48] | select_n2x_8 & (~ IN2[48]) | select_ne_8 & (~ IN2[49])  );
    wire logic pp_8_50;
    assign pp_8_50 = (select_e_8 & IN2[50] | select_2x_8 & IN2[49] | select_n2x_8 & (~ IN2[49]) | select_ne_8 & (~ IN2[50])  );
    wire logic pp_8_51;
    assign pp_8_51 = (select_e_8 & IN2[51] | select_2x_8 & IN2[50] | select_n2x_8 & (~ IN2[50]) | select_ne_8 & (~ IN2[51])  );
    wire logic pp_8_52;
    assign pp_8_52 = (select_e_8 & IN2[52] | select_2x_8 & IN2[51] | select_n2x_8 & (~ IN2[51]) | select_ne_8 & (~ IN2[52])  );
    wire logic pp_8_53;
    assign pp_8_53 = (select_e_8 & IN2[53] | select_2x_8 & IN2[52] | select_n2x_8 & (~ IN2[52]) | select_ne_8 & (~ IN2[53])  );
    wire logic pp_8_54;
    assign pp_8_54 = (select_e_8 & IN2[54] | select_2x_8 & IN2[53] | select_n2x_8 & (~ IN2[53]) | select_ne_8 & (~ IN2[54])  );
    wire logic pp_8_55;
    assign pp_8_55 = (select_e_8 & IN2[55] | select_2x_8 & IN2[54] | select_n2x_8 & (~ IN2[54]) | select_ne_8 & (~ IN2[55])  );
    wire logic pp_8_56;
    assign pp_8_56 = (select_e_8 & IN2[56] | select_2x_8 & IN2[55] | select_n2x_8 & (~ IN2[55]) | select_ne_8 & (~ IN2[56])  );
    wire logic pp_8_57;
    assign pp_8_57 = (select_e_8 & IN2[57] | select_2x_8 & IN2[56] | select_n2x_8 & (~ IN2[56]) | select_ne_8 & (~ IN2[57])  );
    wire logic pp_8_58;
    assign pp_8_58 = (select_e_8 & IN2[58] | select_2x_8 & IN2[57] | select_n2x_8 & (~ IN2[57]) | select_ne_8 & (~ IN2[58])  );
    wire logic pp_8_59;
    assign pp_8_59 = (select_e_8 & IN2[59] | select_2x_8 & IN2[58] | select_n2x_8 & (~ IN2[58]) | select_ne_8 & (~ IN2[59])  );
    wire logic pp_8_60;
    assign pp_8_60 = (select_e_8 & IN2[60] | select_2x_8 & IN2[59] | select_n2x_8 & (~ IN2[59]) | select_ne_8 & (~ IN2[60])  );
    wire logic pp_8_61;
    assign pp_8_61 = (select_e_8 & IN2[61] | select_2x_8 & IN2[60] | select_n2x_8 & (~ IN2[60]) | select_ne_8 & (~ IN2[61])  );
    wire logic pp_8_62;
    assign pp_8_62 = (select_e_8 & IN2[62] | select_2x_8 & IN2[61] | select_n2x_8 & (~ IN2[61]) | select_ne_8 & (~ IN2[62])  );
    wire logic pp_8_63;
    assign pp_8_63 = (select_e_8 & IN2[63] | select_2x_8 & IN2[62] | select_n2x_8 & (~ IN2[62]) | select_ne_8 & (~ IN2[63])  );
    wire logic pp_8_64;
    assign pp_8_64 = (select_e_8 & IN2[63] | select_2x_8 & IN2[63] | select_n2x_8 & (~ IN2[63]) | select_ne_8 & (~ IN2[63])  );
    wire logic pp_8_65;
    assign pp_8_65 = ~ (select_e_8 & IN2[63] | select_2x_8 & IN2[63] | select_n2x_8 & (~ IN2[63]) | select_ne_8 & (~ IN2[63])  );
    assign tcomp8 = select_ne_8 | select_n2x_8;
    
    // Signed Booth Radix-4 Partial Products Row 10
    wire logic select_e_9, select_ne_9, select_2x_9, tcomp9, select_n2x_9;
    assign select_e_9 = ((~ IN1[19]) & (IN1[18] ^ IN1[17]));
    assign select_ne_9 = IN1[19] &  (IN1[18] ^ IN1[17]);
    assign select_2x_9 = (~ IN1[19]) & IN1[18] & IN1[17];
    assign select_n2x_9 = IN1[19] & (~ IN1[18]) & (~ IN1[17]);
    wire logic pp_9_0;
    assign pp_9_0 = (select_e_9 & IN2[0] | select_2x_9 & 1'b0 | select_n2x_9 & 1'b1 | select_ne_9 & (~ IN2[0])  );
    wire logic pp_9_1;
    assign pp_9_1 = (select_e_9 & IN2[1] | select_2x_9 & IN2[0] | select_n2x_9 & (~ IN2[0]) | select_ne_9 & (~ IN2[1])  );
    wire logic pp_9_2;
    assign pp_9_2 = (select_e_9 & IN2[2] | select_2x_9 & IN2[1] | select_n2x_9 & (~ IN2[1]) | select_ne_9 & (~ IN2[2])  );
    wire logic pp_9_3;
    assign pp_9_3 = (select_e_9 & IN2[3] | select_2x_9 & IN2[2] | select_n2x_9 & (~ IN2[2]) | select_ne_9 & (~ IN2[3])  );
    wire logic pp_9_4;
    assign pp_9_4 = (select_e_9 & IN2[4] | select_2x_9 & IN2[3] | select_n2x_9 & (~ IN2[3]) | select_ne_9 & (~ IN2[4])  );
    wire logic pp_9_5;
    assign pp_9_5 = (select_e_9 & IN2[5] | select_2x_9 & IN2[4] | select_n2x_9 & (~ IN2[4]) | select_ne_9 & (~ IN2[5])  );
    wire logic pp_9_6;
    assign pp_9_6 = (select_e_9 & IN2[6] | select_2x_9 & IN2[5] | select_n2x_9 & (~ IN2[5]) | select_ne_9 & (~ IN2[6])  );
    wire logic pp_9_7;
    assign pp_9_7 = (select_e_9 & IN2[7] | select_2x_9 & IN2[6] | select_n2x_9 & (~ IN2[6]) | select_ne_9 & (~ IN2[7])  );
    wire logic pp_9_8;
    assign pp_9_8 = (select_e_9 & IN2[8] | select_2x_9 & IN2[7] | select_n2x_9 & (~ IN2[7]) | select_ne_9 & (~ IN2[8])  );
    wire logic pp_9_9;
    assign pp_9_9 = (select_e_9 & IN2[9] | select_2x_9 & IN2[8] | select_n2x_9 & (~ IN2[8]) | select_ne_9 & (~ IN2[9])  );
    wire logic pp_9_10;
    assign pp_9_10 = (select_e_9 & IN2[10] | select_2x_9 & IN2[9] | select_n2x_9 & (~ IN2[9]) | select_ne_9 & (~ IN2[10])  );
    wire logic pp_9_11;
    assign pp_9_11 = (select_e_9 & IN2[11] | select_2x_9 & IN2[10] | select_n2x_9 & (~ IN2[10]) | select_ne_9 & (~ IN2[11])  );
    wire logic pp_9_12;
    assign pp_9_12 = (select_e_9 & IN2[12] | select_2x_9 & IN2[11] | select_n2x_9 & (~ IN2[11]) | select_ne_9 & (~ IN2[12])  );
    wire logic pp_9_13;
    assign pp_9_13 = (select_e_9 & IN2[13] | select_2x_9 & IN2[12] | select_n2x_9 & (~ IN2[12]) | select_ne_9 & (~ IN2[13])  );
    wire logic pp_9_14;
    assign pp_9_14 = (select_e_9 & IN2[14] | select_2x_9 & IN2[13] | select_n2x_9 & (~ IN2[13]) | select_ne_9 & (~ IN2[14])  );
    wire logic pp_9_15;
    assign pp_9_15 = (select_e_9 & IN2[15] | select_2x_9 & IN2[14] | select_n2x_9 & (~ IN2[14]) | select_ne_9 & (~ IN2[15])  );
    wire logic pp_9_16;
    assign pp_9_16 = (select_e_9 & IN2[16] | select_2x_9 & IN2[15] | select_n2x_9 & (~ IN2[15]) | select_ne_9 & (~ IN2[16])  );
    wire logic pp_9_17;
    assign pp_9_17 = (select_e_9 & IN2[17] | select_2x_9 & IN2[16] | select_n2x_9 & (~ IN2[16]) | select_ne_9 & (~ IN2[17])  );
    wire logic pp_9_18;
    assign pp_9_18 = (select_e_9 & IN2[18] | select_2x_9 & IN2[17] | select_n2x_9 & (~ IN2[17]) | select_ne_9 & (~ IN2[18])  );
    wire logic pp_9_19;
    assign pp_9_19 = (select_e_9 & IN2[19] | select_2x_9 & IN2[18] | select_n2x_9 & (~ IN2[18]) | select_ne_9 & (~ IN2[19])  );
    wire logic pp_9_20;
    assign pp_9_20 = (select_e_9 & IN2[20] | select_2x_9 & IN2[19] | select_n2x_9 & (~ IN2[19]) | select_ne_9 & (~ IN2[20])  );
    wire logic pp_9_21;
    assign pp_9_21 = (select_e_9 & IN2[21] | select_2x_9 & IN2[20] | select_n2x_9 & (~ IN2[20]) | select_ne_9 & (~ IN2[21])  );
    wire logic pp_9_22;
    assign pp_9_22 = (select_e_9 & IN2[22] | select_2x_9 & IN2[21] | select_n2x_9 & (~ IN2[21]) | select_ne_9 & (~ IN2[22])  );
    wire logic pp_9_23;
    assign pp_9_23 = (select_e_9 & IN2[23] | select_2x_9 & IN2[22] | select_n2x_9 & (~ IN2[22]) | select_ne_9 & (~ IN2[23])  );
    wire logic pp_9_24;
    assign pp_9_24 = (select_e_9 & IN2[24] | select_2x_9 & IN2[23] | select_n2x_9 & (~ IN2[23]) | select_ne_9 & (~ IN2[24])  );
    wire logic pp_9_25;
    assign pp_9_25 = (select_e_9 & IN2[25] | select_2x_9 & IN2[24] | select_n2x_9 & (~ IN2[24]) | select_ne_9 & (~ IN2[25])  );
    wire logic pp_9_26;
    assign pp_9_26 = (select_e_9 & IN2[26] | select_2x_9 & IN2[25] | select_n2x_9 & (~ IN2[25]) | select_ne_9 & (~ IN2[26])  );
    wire logic pp_9_27;
    assign pp_9_27 = (select_e_9 & IN2[27] | select_2x_9 & IN2[26] | select_n2x_9 & (~ IN2[26]) | select_ne_9 & (~ IN2[27])  );
    wire logic pp_9_28;
    assign pp_9_28 = (select_e_9 & IN2[28] | select_2x_9 & IN2[27] | select_n2x_9 & (~ IN2[27]) | select_ne_9 & (~ IN2[28])  );
    wire logic pp_9_29;
    assign pp_9_29 = (select_e_9 & IN2[29] | select_2x_9 & IN2[28] | select_n2x_9 & (~ IN2[28]) | select_ne_9 & (~ IN2[29])  );
    wire logic pp_9_30;
    assign pp_9_30 = (select_e_9 & IN2[30] | select_2x_9 & IN2[29] | select_n2x_9 & (~ IN2[29]) | select_ne_9 & (~ IN2[30])  );
    wire logic pp_9_31;
    assign pp_9_31 = (select_e_9 & IN2[31] | select_2x_9 & IN2[30] | select_n2x_9 & (~ IN2[30]) | select_ne_9 & (~ IN2[31])  );
    wire logic pp_9_32;
    assign pp_9_32 = (select_e_9 & IN2[32] | select_2x_9 & IN2[31] | select_n2x_9 & (~ IN2[31]) | select_ne_9 & (~ IN2[32])  );
    wire logic pp_9_33;
    assign pp_9_33 = (select_e_9 & IN2[33] | select_2x_9 & IN2[32] | select_n2x_9 & (~ IN2[32]) | select_ne_9 & (~ IN2[33])  );
    wire logic pp_9_34;
    assign pp_9_34 = (select_e_9 & IN2[34] | select_2x_9 & IN2[33] | select_n2x_9 & (~ IN2[33]) | select_ne_9 & (~ IN2[34])  );
    wire logic pp_9_35;
    assign pp_9_35 = (select_e_9 & IN2[35] | select_2x_9 & IN2[34] | select_n2x_9 & (~ IN2[34]) | select_ne_9 & (~ IN2[35])  );
    wire logic pp_9_36;
    assign pp_9_36 = (select_e_9 & IN2[36] | select_2x_9 & IN2[35] | select_n2x_9 & (~ IN2[35]) | select_ne_9 & (~ IN2[36])  );
    wire logic pp_9_37;
    assign pp_9_37 = (select_e_9 & IN2[37] | select_2x_9 & IN2[36] | select_n2x_9 & (~ IN2[36]) | select_ne_9 & (~ IN2[37])  );
    wire logic pp_9_38;
    assign pp_9_38 = (select_e_9 & IN2[38] | select_2x_9 & IN2[37] | select_n2x_9 & (~ IN2[37]) | select_ne_9 & (~ IN2[38])  );
    wire logic pp_9_39;
    assign pp_9_39 = (select_e_9 & IN2[39] | select_2x_9 & IN2[38] | select_n2x_9 & (~ IN2[38]) | select_ne_9 & (~ IN2[39])  );
    wire logic pp_9_40;
    assign pp_9_40 = (select_e_9 & IN2[40] | select_2x_9 & IN2[39] | select_n2x_9 & (~ IN2[39]) | select_ne_9 & (~ IN2[40])  );
    wire logic pp_9_41;
    assign pp_9_41 = (select_e_9 & IN2[41] | select_2x_9 & IN2[40] | select_n2x_9 & (~ IN2[40]) | select_ne_9 & (~ IN2[41])  );
    wire logic pp_9_42;
    assign pp_9_42 = (select_e_9 & IN2[42] | select_2x_9 & IN2[41] | select_n2x_9 & (~ IN2[41]) | select_ne_9 & (~ IN2[42])  );
    wire logic pp_9_43;
    assign pp_9_43 = (select_e_9 & IN2[43] | select_2x_9 & IN2[42] | select_n2x_9 & (~ IN2[42]) | select_ne_9 & (~ IN2[43])  );
    wire logic pp_9_44;
    assign pp_9_44 = (select_e_9 & IN2[44] | select_2x_9 & IN2[43] | select_n2x_9 & (~ IN2[43]) | select_ne_9 & (~ IN2[44])  );
    wire logic pp_9_45;
    assign pp_9_45 = (select_e_9 & IN2[45] | select_2x_9 & IN2[44] | select_n2x_9 & (~ IN2[44]) | select_ne_9 & (~ IN2[45])  );
    wire logic pp_9_46;
    assign pp_9_46 = (select_e_9 & IN2[46] | select_2x_9 & IN2[45] | select_n2x_9 & (~ IN2[45]) | select_ne_9 & (~ IN2[46])  );
    wire logic pp_9_47;
    assign pp_9_47 = (select_e_9 & IN2[47] | select_2x_9 & IN2[46] | select_n2x_9 & (~ IN2[46]) | select_ne_9 & (~ IN2[47])  );
    wire logic pp_9_48;
    assign pp_9_48 = (select_e_9 & IN2[48] | select_2x_9 & IN2[47] | select_n2x_9 & (~ IN2[47]) | select_ne_9 & (~ IN2[48])  );
    wire logic pp_9_49;
    assign pp_9_49 = (select_e_9 & IN2[49] | select_2x_9 & IN2[48] | select_n2x_9 & (~ IN2[48]) | select_ne_9 & (~ IN2[49])  );
    wire logic pp_9_50;
    assign pp_9_50 = (select_e_9 & IN2[50] | select_2x_9 & IN2[49] | select_n2x_9 & (~ IN2[49]) | select_ne_9 & (~ IN2[50])  );
    wire logic pp_9_51;
    assign pp_9_51 = (select_e_9 & IN2[51] | select_2x_9 & IN2[50] | select_n2x_9 & (~ IN2[50]) | select_ne_9 & (~ IN2[51])  );
    wire logic pp_9_52;
    assign pp_9_52 = (select_e_9 & IN2[52] | select_2x_9 & IN2[51] | select_n2x_9 & (~ IN2[51]) | select_ne_9 & (~ IN2[52])  );
    wire logic pp_9_53;
    assign pp_9_53 = (select_e_9 & IN2[53] | select_2x_9 & IN2[52] | select_n2x_9 & (~ IN2[52]) | select_ne_9 & (~ IN2[53])  );
    wire logic pp_9_54;
    assign pp_9_54 = (select_e_9 & IN2[54] | select_2x_9 & IN2[53] | select_n2x_9 & (~ IN2[53]) | select_ne_9 & (~ IN2[54])  );
    wire logic pp_9_55;
    assign pp_9_55 = (select_e_9 & IN2[55] | select_2x_9 & IN2[54] | select_n2x_9 & (~ IN2[54]) | select_ne_9 & (~ IN2[55])  );
    wire logic pp_9_56;
    assign pp_9_56 = (select_e_9 & IN2[56] | select_2x_9 & IN2[55] | select_n2x_9 & (~ IN2[55]) | select_ne_9 & (~ IN2[56])  );
    wire logic pp_9_57;
    assign pp_9_57 = (select_e_9 & IN2[57] | select_2x_9 & IN2[56] | select_n2x_9 & (~ IN2[56]) | select_ne_9 & (~ IN2[57])  );
    wire logic pp_9_58;
    assign pp_9_58 = (select_e_9 & IN2[58] | select_2x_9 & IN2[57] | select_n2x_9 & (~ IN2[57]) | select_ne_9 & (~ IN2[58])  );
    wire logic pp_9_59;
    assign pp_9_59 = (select_e_9 & IN2[59] | select_2x_9 & IN2[58] | select_n2x_9 & (~ IN2[58]) | select_ne_9 & (~ IN2[59])  );
    wire logic pp_9_60;
    assign pp_9_60 = (select_e_9 & IN2[60] | select_2x_9 & IN2[59] | select_n2x_9 & (~ IN2[59]) | select_ne_9 & (~ IN2[60])  );
    wire logic pp_9_61;
    assign pp_9_61 = (select_e_9 & IN2[61] | select_2x_9 & IN2[60] | select_n2x_9 & (~ IN2[60]) | select_ne_9 & (~ IN2[61])  );
    wire logic pp_9_62;
    assign pp_9_62 = (select_e_9 & IN2[62] | select_2x_9 & IN2[61] | select_n2x_9 & (~ IN2[61]) | select_ne_9 & (~ IN2[62])  );
    wire logic pp_9_63;
    assign pp_9_63 = (select_e_9 & IN2[63] | select_2x_9 & IN2[62] | select_n2x_9 & (~ IN2[62]) | select_ne_9 & (~ IN2[63])  );
    wire logic pp_9_64;
    assign pp_9_64 = (select_e_9 & IN2[63] | select_2x_9 & IN2[63] | select_n2x_9 & (~ IN2[63]) | select_ne_9 & (~ IN2[63])  );
    wire logic pp_9_65;
    assign pp_9_65 = ~ (select_e_9 & IN2[63] | select_2x_9 & IN2[63] | select_n2x_9 & (~ IN2[63]) | select_ne_9 & (~ IN2[63])  );
    assign tcomp9 = select_ne_9 | select_n2x_9;
    
    // Signed Booth Radix-4 Partial Products Row 11
    wire logic select_e_10, select_ne_10, select_2x_10, tcomp10, select_n2x_10;
    assign select_e_10 = ((~ IN1[21]) & (IN1[20] ^ IN1[19]));
    assign select_ne_10 = IN1[21] &  (IN1[20] ^ IN1[19]);
    assign select_2x_10 = (~ IN1[21]) & IN1[20] & IN1[19];
    assign select_n2x_10 = IN1[21] & (~ IN1[20]) & (~ IN1[19]);
    wire logic pp_10_0;
    assign pp_10_0 = (select_e_10 & IN2[0] | select_2x_10 & 1'b0 | select_n2x_10 & 1'b1 | select_ne_10 & (~ IN2[0])  );
    wire logic pp_10_1;
    assign pp_10_1 = (select_e_10 & IN2[1] | select_2x_10 & IN2[0] | select_n2x_10 & (~ IN2[0]) | select_ne_10 & (~ IN2[1])  );
    wire logic pp_10_2;
    assign pp_10_2 = (select_e_10 & IN2[2] | select_2x_10 & IN2[1] | select_n2x_10 & (~ IN2[1]) | select_ne_10 & (~ IN2[2])  );
    wire logic pp_10_3;
    assign pp_10_3 = (select_e_10 & IN2[3] | select_2x_10 & IN2[2] | select_n2x_10 & (~ IN2[2]) | select_ne_10 & (~ IN2[3])  );
    wire logic pp_10_4;
    assign pp_10_4 = (select_e_10 & IN2[4] | select_2x_10 & IN2[3] | select_n2x_10 & (~ IN2[3]) | select_ne_10 & (~ IN2[4])  );
    wire logic pp_10_5;
    assign pp_10_5 = (select_e_10 & IN2[5] | select_2x_10 & IN2[4] | select_n2x_10 & (~ IN2[4]) | select_ne_10 & (~ IN2[5])  );
    wire logic pp_10_6;
    assign pp_10_6 = (select_e_10 & IN2[6] | select_2x_10 & IN2[5] | select_n2x_10 & (~ IN2[5]) | select_ne_10 & (~ IN2[6])  );
    wire logic pp_10_7;
    assign pp_10_7 = (select_e_10 & IN2[7] | select_2x_10 & IN2[6] | select_n2x_10 & (~ IN2[6]) | select_ne_10 & (~ IN2[7])  );
    wire logic pp_10_8;
    assign pp_10_8 = (select_e_10 & IN2[8] | select_2x_10 & IN2[7] | select_n2x_10 & (~ IN2[7]) | select_ne_10 & (~ IN2[8])  );
    wire logic pp_10_9;
    assign pp_10_9 = (select_e_10 & IN2[9] | select_2x_10 & IN2[8] | select_n2x_10 & (~ IN2[8]) | select_ne_10 & (~ IN2[9])  );
    wire logic pp_10_10;
    assign pp_10_10 = (select_e_10 & IN2[10] | select_2x_10 & IN2[9] | select_n2x_10 & (~ IN2[9]) | select_ne_10 & (~ IN2[10])  );
    wire logic pp_10_11;
    assign pp_10_11 = (select_e_10 & IN2[11] | select_2x_10 & IN2[10] | select_n2x_10 & (~ IN2[10]) | select_ne_10 & (~ IN2[11])  );
    wire logic pp_10_12;
    assign pp_10_12 = (select_e_10 & IN2[12] | select_2x_10 & IN2[11] | select_n2x_10 & (~ IN2[11]) | select_ne_10 & (~ IN2[12])  );
    wire logic pp_10_13;
    assign pp_10_13 = (select_e_10 & IN2[13] | select_2x_10 & IN2[12] | select_n2x_10 & (~ IN2[12]) | select_ne_10 & (~ IN2[13])  );
    wire logic pp_10_14;
    assign pp_10_14 = (select_e_10 & IN2[14] | select_2x_10 & IN2[13] | select_n2x_10 & (~ IN2[13]) | select_ne_10 & (~ IN2[14])  );
    wire logic pp_10_15;
    assign pp_10_15 = (select_e_10 & IN2[15] | select_2x_10 & IN2[14] | select_n2x_10 & (~ IN2[14]) | select_ne_10 & (~ IN2[15])  );
    wire logic pp_10_16;
    assign pp_10_16 = (select_e_10 & IN2[16] | select_2x_10 & IN2[15] | select_n2x_10 & (~ IN2[15]) | select_ne_10 & (~ IN2[16])  );
    wire logic pp_10_17;
    assign pp_10_17 = (select_e_10 & IN2[17] | select_2x_10 & IN2[16] | select_n2x_10 & (~ IN2[16]) | select_ne_10 & (~ IN2[17])  );
    wire logic pp_10_18;
    assign pp_10_18 = (select_e_10 & IN2[18] | select_2x_10 & IN2[17] | select_n2x_10 & (~ IN2[17]) | select_ne_10 & (~ IN2[18])  );
    wire logic pp_10_19;
    assign pp_10_19 = (select_e_10 & IN2[19] | select_2x_10 & IN2[18] | select_n2x_10 & (~ IN2[18]) | select_ne_10 & (~ IN2[19])  );
    wire logic pp_10_20;
    assign pp_10_20 = (select_e_10 & IN2[20] | select_2x_10 & IN2[19] | select_n2x_10 & (~ IN2[19]) | select_ne_10 & (~ IN2[20])  );
    wire logic pp_10_21;
    assign pp_10_21 = (select_e_10 & IN2[21] | select_2x_10 & IN2[20] | select_n2x_10 & (~ IN2[20]) | select_ne_10 & (~ IN2[21])  );
    wire logic pp_10_22;
    assign pp_10_22 = (select_e_10 & IN2[22] | select_2x_10 & IN2[21] | select_n2x_10 & (~ IN2[21]) | select_ne_10 & (~ IN2[22])  );
    wire logic pp_10_23;
    assign pp_10_23 = (select_e_10 & IN2[23] | select_2x_10 & IN2[22] | select_n2x_10 & (~ IN2[22]) | select_ne_10 & (~ IN2[23])  );
    wire logic pp_10_24;
    assign pp_10_24 = (select_e_10 & IN2[24] | select_2x_10 & IN2[23] | select_n2x_10 & (~ IN2[23]) | select_ne_10 & (~ IN2[24])  );
    wire logic pp_10_25;
    assign pp_10_25 = (select_e_10 & IN2[25] | select_2x_10 & IN2[24] | select_n2x_10 & (~ IN2[24]) | select_ne_10 & (~ IN2[25])  );
    wire logic pp_10_26;
    assign pp_10_26 = (select_e_10 & IN2[26] | select_2x_10 & IN2[25] | select_n2x_10 & (~ IN2[25]) | select_ne_10 & (~ IN2[26])  );
    wire logic pp_10_27;
    assign pp_10_27 = (select_e_10 & IN2[27] | select_2x_10 & IN2[26] | select_n2x_10 & (~ IN2[26]) | select_ne_10 & (~ IN2[27])  );
    wire logic pp_10_28;
    assign pp_10_28 = (select_e_10 & IN2[28] | select_2x_10 & IN2[27] | select_n2x_10 & (~ IN2[27]) | select_ne_10 & (~ IN2[28])  );
    wire logic pp_10_29;
    assign pp_10_29 = (select_e_10 & IN2[29] | select_2x_10 & IN2[28] | select_n2x_10 & (~ IN2[28]) | select_ne_10 & (~ IN2[29])  );
    wire logic pp_10_30;
    assign pp_10_30 = (select_e_10 & IN2[30] | select_2x_10 & IN2[29] | select_n2x_10 & (~ IN2[29]) | select_ne_10 & (~ IN2[30])  );
    wire logic pp_10_31;
    assign pp_10_31 = (select_e_10 & IN2[31] | select_2x_10 & IN2[30] | select_n2x_10 & (~ IN2[30]) | select_ne_10 & (~ IN2[31])  );
    wire logic pp_10_32;
    assign pp_10_32 = (select_e_10 & IN2[32] | select_2x_10 & IN2[31] | select_n2x_10 & (~ IN2[31]) | select_ne_10 & (~ IN2[32])  );
    wire logic pp_10_33;
    assign pp_10_33 = (select_e_10 & IN2[33] | select_2x_10 & IN2[32] | select_n2x_10 & (~ IN2[32]) | select_ne_10 & (~ IN2[33])  );
    wire logic pp_10_34;
    assign pp_10_34 = (select_e_10 & IN2[34] | select_2x_10 & IN2[33] | select_n2x_10 & (~ IN2[33]) | select_ne_10 & (~ IN2[34])  );
    wire logic pp_10_35;
    assign pp_10_35 = (select_e_10 & IN2[35] | select_2x_10 & IN2[34] | select_n2x_10 & (~ IN2[34]) | select_ne_10 & (~ IN2[35])  );
    wire logic pp_10_36;
    assign pp_10_36 = (select_e_10 & IN2[36] | select_2x_10 & IN2[35] | select_n2x_10 & (~ IN2[35]) | select_ne_10 & (~ IN2[36])  );
    wire logic pp_10_37;
    assign pp_10_37 = (select_e_10 & IN2[37] | select_2x_10 & IN2[36] | select_n2x_10 & (~ IN2[36]) | select_ne_10 & (~ IN2[37])  );
    wire logic pp_10_38;
    assign pp_10_38 = (select_e_10 & IN2[38] | select_2x_10 & IN2[37] | select_n2x_10 & (~ IN2[37]) | select_ne_10 & (~ IN2[38])  );
    wire logic pp_10_39;
    assign pp_10_39 = (select_e_10 & IN2[39] | select_2x_10 & IN2[38] | select_n2x_10 & (~ IN2[38]) | select_ne_10 & (~ IN2[39])  );
    wire logic pp_10_40;
    assign pp_10_40 = (select_e_10 & IN2[40] | select_2x_10 & IN2[39] | select_n2x_10 & (~ IN2[39]) | select_ne_10 & (~ IN2[40])  );
    wire logic pp_10_41;
    assign pp_10_41 = (select_e_10 & IN2[41] | select_2x_10 & IN2[40] | select_n2x_10 & (~ IN2[40]) | select_ne_10 & (~ IN2[41])  );
    wire logic pp_10_42;
    assign pp_10_42 = (select_e_10 & IN2[42] | select_2x_10 & IN2[41] | select_n2x_10 & (~ IN2[41]) | select_ne_10 & (~ IN2[42])  );
    wire logic pp_10_43;
    assign pp_10_43 = (select_e_10 & IN2[43] | select_2x_10 & IN2[42] | select_n2x_10 & (~ IN2[42]) | select_ne_10 & (~ IN2[43])  );
    wire logic pp_10_44;
    assign pp_10_44 = (select_e_10 & IN2[44] | select_2x_10 & IN2[43] | select_n2x_10 & (~ IN2[43]) | select_ne_10 & (~ IN2[44])  );
    wire logic pp_10_45;
    assign pp_10_45 = (select_e_10 & IN2[45] | select_2x_10 & IN2[44] | select_n2x_10 & (~ IN2[44]) | select_ne_10 & (~ IN2[45])  );
    wire logic pp_10_46;
    assign pp_10_46 = (select_e_10 & IN2[46] | select_2x_10 & IN2[45] | select_n2x_10 & (~ IN2[45]) | select_ne_10 & (~ IN2[46])  );
    wire logic pp_10_47;
    assign pp_10_47 = (select_e_10 & IN2[47] | select_2x_10 & IN2[46] | select_n2x_10 & (~ IN2[46]) | select_ne_10 & (~ IN2[47])  );
    wire logic pp_10_48;
    assign pp_10_48 = (select_e_10 & IN2[48] | select_2x_10 & IN2[47] | select_n2x_10 & (~ IN2[47]) | select_ne_10 & (~ IN2[48])  );
    wire logic pp_10_49;
    assign pp_10_49 = (select_e_10 & IN2[49] | select_2x_10 & IN2[48] | select_n2x_10 & (~ IN2[48]) | select_ne_10 & (~ IN2[49])  );
    wire logic pp_10_50;
    assign pp_10_50 = (select_e_10 & IN2[50] | select_2x_10 & IN2[49] | select_n2x_10 & (~ IN2[49]) | select_ne_10 & (~ IN2[50])  );
    wire logic pp_10_51;
    assign pp_10_51 = (select_e_10 & IN2[51] | select_2x_10 & IN2[50] | select_n2x_10 & (~ IN2[50]) | select_ne_10 & (~ IN2[51])  );
    wire logic pp_10_52;
    assign pp_10_52 = (select_e_10 & IN2[52] | select_2x_10 & IN2[51] | select_n2x_10 & (~ IN2[51]) | select_ne_10 & (~ IN2[52])  );
    wire logic pp_10_53;
    assign pp_10_53 = (select_e_10 & IN2[53] | select_2x_10 & IN2[52] | select_n2x_10 & (~ IN2[52]) | select_ne_10 & (~ IN2[53])  );
    wire logic pp_10_54;
    assign pp_10_54 = (select_e_10 & IN2[54] | select_2x_10 & IN2[53] | select_n2x_10 & (~ IN2[53]) | select_ne_10 & (~ IN2[54])  );
    wire logic pp_10_55;
    assign pp_10_55 = (select_e_10 & IN2[55] | select_2x_10 & IN2[54] | select_n2x_10 & (~ IN2[54]) | select_ne_10 & (~ IN2[55])  );
    wire logic pp_10_56;
    assign pp_10_56 = (select_e_10 & IN2[56] | select_2x_10 & IN2[55] | select_n2x_10 & (~ IN2[55]) | select_ne_10 & (~ IN2[56])  );
    wire logic pp_10_57;
    assign pp_10_57 = (select_e_10 & IN2[57] | select_2x_10 & IN2[56] | select_n2x_10 & (~ IN2[56]) | select_ne_10 & (~ IN2[57])  );
    wire logic pp_10_58;
    assign pp_10_58 = (select_e_10 & IN2[58] | select_2x_10 & IN2[57] | select_n2x_10 & (~ IN2[57]) | select_ne_10 & (~ IN2[58])  );
    wire logic pp_10_59;
    assign pp_10_59 = (select_e_10 & IN2[59] | select_2x_10 & IN2[58] | select_n2x_10 & (~ IN2[58]) | select_ne_10 & (~ IN2[59])  );
    wire logic pp_10_60;
    assign pp_10_60 = (select_e_10 & IN2[60] | select_2x_10 & IN2[59] | select_n2x_10 & (~ IN2[59]) | select_ne_10 & (~ IN2[60])  );
    wire logic pp_10_61;
    assign pp_10_61 = (select_e_10 & IN2[61] | select_2x_10 & IN2[60] | select_n2x_10 & (~ IN2[60]) | select_ne_10 & (~ IN2[61])  );
    wire logic pp_10_62;
    assign pp_10_62 = (select_e_10 & IN2[62] | select_2x_10 & IN2[61] | select_n2x_10 & (~ IN2[61]) | select_ne_10 & (~ IN2[62])  );
    wire logic pp_10_63;
    assign pp_10_63 = (select_e_10 & IN2[63] | select_2x_10 & IN2[62] | select_n2x_10 & (~ IN2[62]) | select_ne_10 & (~ IN2[63])  );
    wire logic pp_10_64;
    assign pp_10_64 = (select_e_10 & IN2[63] | select_2x_10 & IN2[63] | select_n2x_10 & (~ IN2[63]) | select_ne_10 & (~ IN2[63])  );
    wire logic pp_10_65;
    assign pp_10_65 = ~ (select_e_10 & IN2[63] | select_2x_10 & IN2[63] | select_n2x_10 & (~ IN2[63]) | select_ne_10 & (~ IN2[63])  );
    assign tcomp10 = select_ne_10 | select_n2x_10;
    
    // Signed Booth Radix-4 Partial Products Row 12
    wire logic select_e_11, select_ne_11, select_2x_11, tcomp11, select_n2x_11;
    assign select_e_11 = ((~ IN1[23]) & (IN1[22] ^ IN1[21]));
    assign select_ne_11 = IN1[23] &  (IN1[22] ^ IN1[21]);
    assign select_2x_11 = (~ IN1[23]) & IN1[22] & IN1[21];
    assign select_n2x_11 = IN1[23] & (~ IN1[22]) & (~ IN1[21]);
    wire logic pp_11_0;
    assign pp_11_0 = (select_e_11 & IN2[0] | select_2x_11 & 1'b0 | select_n2x_11 & 1'b1 | select_ne_11 & (~ IN2[0])  );
    wire logic pp_11_1;
    assign pp_11_1 = (select_e_11 & IN2[1] | select_2x_11 & IN2[0] | select_n2x_11 & (~ IN2[0]) | select_ne_11 & (~ IN2[1])  );
    wire logic pp_11_2;
    assign pp_11_2 = (select_e_11 & IN2[2] | select_2x_11 & IN2[1] | select_n2x_11 & (~ IN2[1]) | select_ne_11 & (~ IN2[2])  );
    wire logic pp_11_3;
    assign pp_11_3 = (select_e_11 & IN2[3] | select_2x_11 & IN2[2] | select_n2x_11 & (~ IN2[2]) | select_ne_11 & (~ IN2[3])  );
    wire logic pp_11_4;
    assign pp_11_4 = (select_e_11 & IN2[4] | select_2x_11 & IN2[3] | select_n2x_11 & (~ IN2[3]) | select_ne_11 & (~ IN2[4])  );
    wire logic pp_11_5;
    assign pp_11_5 = (select_e_11 & IN2[5] | select_2x_11 & IN2[4] | select_n2x_11 & (~ IN2[4]) | select_ne_11 & (~ IN2[5])  );
    wire logic pp_11_6;
    assign pp_11_6 = (select_e_11 & IN2[6] | select_2x_11 & IN2[5] | select_n2x_11 & (~ IN2[5]) | select_ne_11 & (~ IN2[6])  );
    wire logic pp_11_7;
    assign pp_11_7 = (select_e_11 & IN2[7] | select_2x_11 & IN2[6] | select_n2x_11 & (~ IN2[6]) | select_ne_11 & (~ IN2[7])  );
    wire logic pp_11_8;
    assign pp_11_8 = (select_e_11 & IN2[8] | select_2x_11 & IN2[7] | select_n2x_11 & (~ IN2[7]) | select_ne_11 & (~ IN2[8])  );
    wire logic pp_11_9;
    assign pp_11_9 = (select_e_11 & IN2[9] | select_2x_11 & IN2[8] | select_n2x_11 & (~ IN2[8]) | select_ne_11 & (~ IN2[9])  );
    wire logic pp_11_10;
    assign pp_11_10 = (select_e_11 & IN2[10] | select_2x_11 & IN2[9] | select_n2x_11 & (~ IN2[9]) | select_ne_11 & (~ IN2[10])  );
    wire logic pp_11_11;
    assign pp_11_11 = (select_e_11 & IN2[11] | select_2x_11 & IN2[10] | select_n2x_11 & (~ IN2[10]) | select_ne_11 & (~ IN2[11])  );
    wire logic pp_11_12;
    assign pp_11_12 = (select_e_11 & IN2[12] | select_2x_11 & IN2[11] | select_n2x_11 & (~ IN2[11]) | select_ne_11 & (~ IN2[12])  );
    wire logic pp_11_13;
    assign pp_11_13 = (select_e_11 & IN2[13] | select_2x_11 & IN2[12] | select_n2x_11 & (~ IN2[12]) | select_ne_11 & (~ IN2[13])  );
    wire logic pp_11_14;
    assign pp_11_14 = (select_e_11 & IN2[14] | select_2x_11 & IN2[13] | select_n2x_11 & (~ IN2[13]) | select_ne_11 & (~ IN2[14])  );
    wire logic pp_11_15;
    assign pp_11_15 = (select_e_11 & IN2[15] | select_2x_11 & IN2[14] | select_n2x_11 & (~ IN2[14]) | select_ne_11 & (~ IN2[15])  );
    wire logic pp_11_16;
    assign pp_11_16 = (select_e_11 & IN2[16] | select_2x_11 & IN2[15] | select_n2x_11 & (~ IN2[15]) | select_ne_11 & (~ IN2[16])  );
    wire logic pp_11_17;
    assign pp_11_17 = (select_e_11 & IN2[17] | select_2x_11 & IN2[16] | select_n2x_11 & (~ IN2[16]) | select_ne_11 & (~ IN2[17])  );
    wire logic pp_11_18;
    assign pp_11_18 = (select_e_11 & IN2[18] | select_2x_11 & IN2[17] | select_n2x_11 & (~ IN2[17]) | select_ne_11 & (~ IN2[18])  );
    wire logic pp_11_19;
    assign pp_11_19 = (select_e_11 & IN2[19] | select_2x_11 & IN2[18] | select_n2x_11 & (~ IN2[18]) | select_ne_11 & (~ IN2[19])  );
    wire logic pp_11_20;
    assign pp_11_20 = (select_e_11 & IN2[20] | select_2x_11 & IN2[19] | select_n2x_11 & (~ IN2[19]) | select_ne_11 & (~ IN2[20])  );
    wire logic pp_11_21;
    assign pp_11_21 = (select_e_11 & IN2[21] | select_2x_11 & IN2[20] | select_n2x_11 & (~ IN2[20]) | select_ne_11 & (~ IN2[21])  );
    wire logic pp_11_22;
    assign pp_11_22 = (select_e_11 & IN2[22] | select_2x_11 & IN2[21] | select_n2x_11 & (~ IN2[21]) | select_ne_11 & (~ IN2[22])  );
    wire logic pp_11_23;
    assign pp_11_23 = (select_e_11 & IN2[23] | select_2x_11 & IN2[22] | select_n2x_11 & (~ IN2[22]) | select_ne_11 & (~ IN2[23])  );
    wire logic pp_11_24;
    assign pp_11_24 = (select_e_11 & IN2[24] | select_2x_11 & IN2[23] | select_n2x_11 & (~ IN2[23]) | select_ne_11 & (~ IN2[24])  );
    wire logic pp_11_25;
    assign pp_11_25 = (select_e_11 & IN2[25] | select_2x_11 & IN2[24] | select_n2x_11 & (~ IN2[24]) | select_ne_11 & (~ IN2[25])  );
    wire logic pp_11_26;
    assign pp_11_26 = (select_e_11 & IN2[26] | select_2x_11 & IN2[25] | select_n2x_11 & (~ IN2[25]) | select_ne_11 & (~ IN2[26])  );
    wire logic pp_11_27;
    assign pp_11_27 = (select_e_11 & IN2[27] | select_2x_11 & IN2[26] | select_n2x_11 & (~ IN2[26]) | select_ne_11 & (~ IN2[27])  );
    wire logic pp_11_28;
    assign pp_11_28 = (select_e_11 & IN2[28] | select_2x_11 & IN2[27] | select_n2x_11 & (~ IN2[27]) | select_ne_11 & (~ IN2[28])  );
    wire logic pp_11_29;
    assign pp_11_29 = (select_e_11 & IN2[29] | select_2x_11 & IN2[28] | select_n2x_11 & (~ IN2[28]) | select_ne_11 & (~ IN2[29])  );
    wire logic pp_11_30;
    assign pp_11_30 = (select_e_11 & IN2[30] | select_2x_11 & IN2[29] | select_n2x_11 & (~ IN2[29]) | select_ne_11 & (~ IN2[30])  );
    wire logic pp_11_31;
    assign pp_11_31 = (select_e_11 & IN2[31] | select_2x_11 & IN2[30] | select_n2x_11 & (~ IN2[30]) | select_ne_11 & (~ IN2[31])  );
    wire logic pp_11_32;
    assign pp_11_32 = (select_e_11 & IN2[32] | select_2x_11 & IN2[31] | select_n2x_11 & (~ IN2[31]) | select_ne_11 & (~ IN2[32])  );
    wire logic pp_11_33;
    assign pp_11_33 = (select_e_11 & IN2[33] | select_2x_11 & IN2[32] | select_n2x_11 & (~ IN2[32]) | select_ne_11 & (~ IN2[33])  );
    wire logic pp_11_34;
    assign pp_11_34 = (select_e_11 & IN2[34] | select_2x_11 & IN2[33] | select_n2x_11 & (~ IN2[33]) | select_ne_11 & (~ IN2[34])  );
    wire logic pp_11_35;
    assign pp_11_35 = (select_e_11 & IN2[35] | select_2x_11 & IN2[34] | select_n2x_11 & (~ IN2[34]) | select_ne_11 & (~ IN2[35])  );
    wire logic pp_11_36;
    assign pp_11_36 = (select_e_11 & IN2[36] | select_2x_11 & IN2[35] | select_n2x_11 & (~ IN2[35]) | select_ne_11 & (~ IN2[36])  );
    wire logic pp_11_37;
    assign pp_11_37 = (select_e_11 & IN2[37] | select_2x_11 & IN2[36] | select_n2x_11 & (~ IN2[36]) | select_ne_11 & (~ IN2[37])  );
    wire logic pp_11_38;
    assign pp_11_38 = (select_e_11 & IN2[38] | select_2x_11 & IN2[37] | select_n2x_11 & (~ IN2[37]) | select_ne_11 & (~ IN2[38])  );
    wire logic pp_11_39;
    assign pp_11_39 = (select_e_11 & IN2[39] | select_2x_11 & IN2[38] | select_n2x_11 & (~ IN2[38]) | select_ne_11 & (~ IN2[39])  );
    wire logic pp_11_40;
    assign pp_11_40 = (select_e_11 & IN2[40] | select_2x_11 & IN2[39] | select_n2x_11 & (~ IN2[39]) | select_ne_11 & (~ IN2[40])  );
    wire logic pp_11_41;
    assign pp_11_41 = (select_e_11 & IN2[41] | select_2x_11 & IN2[40] | select_n2x_11 & (~ IN2[40]) | select_ne_11 & (~ IN2[41])  );
    wire logic pp_11_42;
    assign pp_11_42 = (select_e_11 & IN2[42] | select_2x_11 & IN2[41] | select_n2x_11 & (~ IN2[41]) | select_ne_11 & (~ IN2[42])  );
    wire logic pp_11_43;
    assign pp_11_43 = (select_e_11 & IN2[43] | select_2x_11 & IN2[42] | select_n2x_11 & (~ IN2[42]) | select_ne_11 & (~ IN2[43])  );
    wire logic pp_11_44;
    assign pp_11_44 = (select_e_11 & IN2[44] | select_2x_11 & IN2[43] | select_n2x_11 & (~ IN2[43]) | select_ne_11 & (~ IN2[44])  );
    wire logic pp_11_45;
    assign pp_11_45 = (select_e_11 & IN2[45] | select_2x_11 & IN2[44] | select_n2x_11 & (~ IN2[44]) | select_ne_11 & (~ IN2[45])  );
    wire logic pp_11_46;
    assign pp_11_46 = (select_e_11 & IN2[46] | select_2x_11 & IN2[45] | select_n2x_11 & (~ IN2[45]) | select_ne_11 & (~ IN2[46])  );
    wire logic pp_11_47;
    assign pp_11_47 = (select_e_11 & IN2[47] | select_2x_11 & IN2[46] | select_n2x_11 & (~ IN2[46]) | select_ne_11 & (~ IN2[47])  );
    wire logic pp_11_48;
    assign pp_11_48 = (select_e_11 & IN2[48] | select_2x_11 & IN2[47] | select_n2x_11 & (~ IN2[47]) | select_ne_11 & (~ IN2[48])  );
    wire logic pp_11_49;
    assign pp_11_49 = (select_e_11 & IN2[49] | select_2x_11 & IN2[48] | select_n2x_11 & (~ IN2[48]) | select_ne_11 & (~ IN2[49])  );
    wire logic pp_11_50;
    assign pp_11_50 = (select_e_11 & IN2[50] | select_2x_11 & IN2[49] | select_n2x_11 & (~ IN2[49]) | select_ne_11 & (~ IN2[50])  );
    wire logic pp_11_51;
    assign pp_11_51 = (select_e_11 & IN2[51] | select_2x_11 & IN2[50] | select_n2x_11 & (~ IN2[50]) | select_ne_11 & (~ IN2[51])  );
    wire logic pp_11_52;
    assign pp_11_52 = (select_e_11 & IN2[52] | select_2x_11 & IN2[51] | select_n2x_11 & (~ IN2[51]) | select_ne_11 & (~ IN2[52])  );
    wire logic pp_11_53;
    assign pp_11_53 = (select_e_11 & IN2[53] | select_2x_11 & IN2[52] | select_n2x_11 & (~ IN2[52]) | select_ne_11 & (~ IN2[53])  );
    wire logic pp_11_54;
    assign pp_11_54 = (select_e_11 & IN2[54] | select_2x_11 & IN2[53] | select_n2x_11 & (~ IN2[53]) | select_ne_11 & (~ IN2[54])  );
    wire logic pp_11_55;
    assign pp_11_55 = (select_e_11 & IN2[55] | select_2x_11 & IN2[54] | select_n2x_11 & (~ IN2[54]) | select_ne_11 & (~ IN2[55])  );
    wire logic pp_11_56;
    assign pp_11_56 = (select_e_11 & IN2[56] | select_2x_11 & IN2[55] | select_n2x_11 & (~ IN2[55]) | select_ne_11 & (~ IN2[56])  );
    wire logic pp_11_57;
    assign pp_11_57 = (select_e_11 & IN2[57] | select_2x_11 & IN2[56] | select_n2x_11 & (~ IN2[56]) | select_ne_11 & (~ IN2[57])  );
    wire logic pp_11_58;
    assign pp_11_58 = (select_e_11 & IN2[58] | select_2x_11 & IN2[57] | select_n2x_11 & (~ IN2[57]) | select_ne_11 & (~ IN2[58])  );
    wire logic pp_11_59;
    assign pp_11_59 = (select_e_11 & IN2[59] | select_2x_11 & IN2[58] | select_n2x_11 & (~ IN2[58]) | select_ne_11 & (~ IN2[59])  );
    wire logic pp_11_60;
    assign pp_11_60 = (select_e_11 & IN2[60] | select_2x_11 & IN2[59] | select_n2x_11 & (~ IN2[59]) | select_ne_11 & (~ IN2[60])  );
    wire logic pp_11_61;
    assign pp_11_61 = (select_e_11 & IN2[61] | select_2x_11 & IN2[60] | select_n2x_11 & (~ IN2[60]) | select_ne_11 & (~ IN2[61])  );
    wire logic pp_11_62;
    assign pp_11_62 = (select_e_11 & IN2[62] | select_2x_11 & IN2[61] | select_n2x_11 & (~ IN2[61]) | select_ne_11 & (~ IN2[62])  );
    wire logic pp_11_63;
    assign pp_11_63 = (select_e_11 & IN2[63] | select_2x_11 & IN2[62] | select_n2x_11 & (~ IN2[62]) | select_ne_11 & (~ IN2[63])  );
    wire logic pp_11_64;
    assign pp_11_64 = (select_e_11 & IN2[63] | select_2x_11 & IN2[63] | select_n2x_11 & (~ IN2[63]) | select_ne_11 & (~ IN2[63])  );
    wire logic pp_11_65;
    assign pp_11_65 = ~ (select_e_11 & IN2[63] | select_2x_11 & IN2[63] | select_n2x_11 & (~ IN2[63]) | select_ne_11 & (~ IN2[63])  );
    assign tcomp11 = select_ne_11 | select_n2x_11;
    
    // Signed Booth Radix-4 Partial Products Row 13
    wire logic select_e_12, select_ne_12, select_2x_12, tcomp12, select_n2x_12;
    assign select_e_12 = ((~ IN1[25]) & (IN1[24] ^ IN1[23]));
    assign select_ne_12 = IN1[25] &  (IN1[24] ^ IN1[23]);
    assign select_2x_12 = (~ IN1[25]) & IN1[24] & IN1[23];
    assign select_n2x_12 = IN1[25] & (~ IN1[24]) & (~ IN1[23]);
    wire logic pp_12_0;
    assign pp_12_0 = (select_e_12 & IN2[0] | select_2x_12 & 1'b0 | select_n2x_12 & 1'b1 | select_ne_12 & (~ IN2[0])  );
    wire logic pp_12_1;
    assign pp_12_1 = (select_e_12 & IN2[1] | select_2x_12 & IN2[0] | select_n2x_12 & (~ IN2[0]) | select_ne_12 & (~ IN2[1])  );
    wire logic pp_12_2;
    assign pp_12_2 = (select_e_12 & IN2[2] | select_2x_12 & IN2[1] | select_n2x_12 & (~ IN2[1]) | select_ne_12 & (~ IN2[2])  );
    wire logic pp_12_3;
    assign pp_12_3 = (select_e_12 & IN2[3] | select_2x_12 & IN2[2] | select_n2x_12 & (~ IN2[2]) | select_ne_12 & (~ IN2[3])  );
    wire logic pp_12_4;
    assign pp_12_4 = (select_e_12 & IN2[4] | select_2x_12 & IN2[3] | select_n2x_12 & (~ IN2[3]) | select_ne_12 & (~ IN2[4])  );
    wire logic pp_12_5;
    assign pp_12_5 = (select_e_12 & IN2[5] | select_2x_12 & IN2[4] | select_n2x_12 & (~ IN2[4]) | select_ne_12 & (~ IN2[5])  );
    wire logic pp_12_6;
    assign pp_12_6 = (select_e_12 & IN2[6] | select_2x_12 & IN2[5] | select_n2x_12 & (~ IN2[5]) | select_ne_12 & (~ IN2[6])  );
    wire logic pp_12_7;
    assign pp_12_7 = (select_e_12 & IN2[7] | select_2x_12 & IN2[6] | select_n2x_12 & (~ IN2[6]) | select_ne_12 & (~ IN2[7])  );
    wire logic pp_12_8;
    assign pp_12_8 = (select_e_12 & IN2[8] | select_2x_12 & IN2[7] | select_n2x_12 & (~ IN2[7]) | select_ne_12 & (~ IN2[8])  );
    wire logic pp_12_9;
    assign pp_12_9 = (select_e_12 & IN2[9] | select_2x_12 & IN2[8] | select_n2x_12 & (~ IN2[8]) | select_ne_12 & (~ IN2[9])  );
    wire logic pp_12_10;
    assign pp_12_10 = (select_e_12 & IN2[10] | select_2x_12 & IN2[9] | select_n2x_12 & (~ IN2[9]) | select_ne_12 & (~ IN2[10])  );
    wire logic pp_12_11;
    assign pp_12_11 = (select_e_12 & IN2[11] | select_2x_12 & IN2[10] | select_n2x_12 & (~ IN2[10]) | select_ne_12 & (~ IN2[11])  );
    wire logic pp_12_12;
    assign pp_12_12 = (select_e_12 & IN2[12] | select_2x_12 & IN2[11] | select_n2x_12 & (~ IN2[11]) | select_ne_12 & (~ IN2[12])  );
    wire logic pp_12_13;
    assign pp_12_13 = (select_e_12 & IN2[13] | select_2x_12 & IN2[12] | select_n2x_12 & (~ IN2[12]) | select_ne_12 & (~ IN2[13])  );
    wire logic pp_12_14;
    assign pp_12_14 = (select_e_12 & IN2[14] | select_2x_12 & IN2[13] | select_n2x_12 & (~ IN2[13]) | select_ne_12 & (~ IN2[14])  );
    wire logic pp_12_15;
    assign pp_12_15 = (select_e_12 & IN2[15] | select_2x_12 & IN2[14] | select_n2x_12 & (~ IN2[14]) | select_ne_12 & (~ IN2[15])  );
    wire logic pp_12_16;
    assign pp_12_16 = (select_e_12 & IN2[16] | select_2x_12 & IN2[15] | select_n2x_12 & (~ IN2[15]) | select_ne_12 & (~ IN2[16])  );
    wire logic pp_12_17;
    assign pp_12_17 = (select_e_12 & IN2[17] | select_2x_12 & IN2[16] | select_n2x_12 & (~ IN2[16]) | select_ne_12 & (~ IN2[17])  );
    wire logic pp_12_18;
    assign pp_12_18 = (select_e_12 & IN2[18] | select_2x_12 & IN2[17] | select_n2x_12 & (~ IN2[17]) | select_ne_12 & (~ IN2[18])  );
    wire logic pp_12_19;
    assign pp_12_19 = (select_e_12 & IN2[19] | select_2x_12 & IN2[18] | select_n2x_12 & (~ IN2[18]) | select_ne_12 & (~ IN2[19])  );
    wire logic pp_12_20;
    assign pp_12_20 = (select_e_12 & IN2[20] | select_2x_12 & IN2[19] | select_n2x_12 & (~ IN2[19]) | select_ne_12 & (~ IN2[20])  );
    wire logic pp_12_21;
    assign pp_12_21 = (select_e_12 & IN2[21] | select_2x_12 & IN2[20] | select_n2x_12 & (~ IN2[20]) | select_ne_12 & (~ IN2[21])  );
    wire logic pp_12_22;
    assign pp_12_22 = (select_e_12 & IN2[22] | select_2x_12 & IN2[21] | select_n2x_12 & (~ IN2[21]) | select_ne_12 & (~ IN2[22])  );
    wire logic pp_12_23;
    assign pp_12_23 = (select_e_12 & IN2[23] | select_2x_12 & IN2[22] | select_n2x_12 & (~ IN2[22]) | select_ne_12 & (~ IN2[23])  );
    wire logic pp_12_24;
    assign pp_12_24 = (select_e_12 & IN2[24] | select_2x_12 & IN2[23] | select_n2x_12 & (~ IN2[23]) | select_ne_12 & (~ IN2[24])  );
    wire logic pp_12_25;
    assign pp_12_25 = (select_e_12 & IN2[25] | select_2x_12 & IN2[24] | select_n2x_12 & (~ IN2[24]) | select_ne_12 & (~ IN2[25])  );
    wire logic pp_12_26;
    assign pp_12_26 = (select_e_12 & IN2[26] | select_2x_12 & IN2[25] | select_n2x_12 & (~ IN2[25]) | select_ne_12 & (~ IN2[26])  );
    wire logic pp_12_27;
    assign pp_12_27 = (select_e_12 & IN2[27] | select_2x_12 & IN2[26] | select_n2x_12 & (~ IN2[26]) | select_ne_12 & (~ IN2[27])  );
    wire logic pp_12_28;
    assign pp_12_28 = (select_e_12 & IN2[28] | select_2x_12 & IN2[27] | select_n2x_12 & (~ IN2[27]) | select_ne_12 & (~ IN2[28])  );
    wire logic pp_12_29;
    assign pp_12_29 = (select_e_12 & IN2[29] | select_2x_12 & IN2[28] | select_n2x_12 & (~ IN2[28]) | select_ne_12 & (~ IN2[29])  );
    wire logic pp_12_30;
    assign pp_12_30 = (select_e_12 & IN2[30] | select_2x_12 & IN2[29] | select_n2x_12 & (~ IN2[29]) | select_ne_12 & (~ IN2[30])  );
    wire logic pp_12_31;
    assign pp_12_31 = (select_e_12 & IN2[31] | select_2x_12 & IN2[30] | select_n2x_12 & (~ IN2[30]) | select_ne_12 & (~ IN2[31])  );
    wire logic pp_12_32;
    assign pp_12_32 = (select_e_12 & IN2[32] | select_2x_12 & IN2[31] | select_n2x_12 & (~ IN2[31]) | select_ne_12 & (~ IN2[32])  );
    wire logic pp_12_33;
    assign pp_12_33 = (select_e_12 & IN2[33] | select_2x_12 & IN2[32] | select_n2x_12 & (~ IN2[32]) | select_ne_12 & (~ IN2[33])  );
    wire logic pp_12_34;
    assign pp_12_34 = (select_e_12 & IN2[34] | select_2x_12 & IN2[33] | select_n2x_12 & (~ IN2[33]) | select_ne_12 & (~ IN2[34])  );
    wire logic pp_12_35;
    assign pp_12_35 = (select_e_12 & IN2[35] | select_2x_12 & IN2[34] | select_n2x_12 & (~ IN2[34]) | select_ne_12 & (~ IN2[35])  );
    wire logic pp_12_36;
    assign pp_12_36 = (select_e_12 & IN2[36] | select_2x_12 & IN2[35] | select_n2x_12 & (~ IN2[35]) | select_ne_12 & (~ IN2[36])  );
    wire logic pp_12_37;
    assign pp_12_37 = (select_e_12 & IN2[37] | select_2x_12 & IN2[36] | select_n2x_12 & (~ IN2[36]) | select_ne_12 & (~ IN2[37])  );
    wire logic pp_12_38;
    assign pp_12_38 = (select_e_12 & IN2[38] | select_2x_12 & IN2[37] | select_n2x_12 & (~ IN2[37]) | select_ne_12 & (~ IN2[38])  );
    wire logic pp_12_39;
    assign pp_12_39 = (select_e_12 & IN2[39] | select_2x_12 & IN2[38] | select_n2x_12 & (~ IN2[38]) | select_ne_12 & (~ IN2[39])  );
    wire logic pp_12_40;
    assign pp_12_40 = (select_e_12 & IN2[40] | select_2x_12 & IN2[39] | select_n2x_12 & (~ IN2[39]) | select_ne_12 & (~ IN2[40])  );
    wire logic pp_12_41;
    assign pp_12_41 = (select_e_12 & IN2[41] | select_2x_12 & IN2[40] | select_n2x_12 & (~ IN2[40]) | select_ne_12 & (~ IN2[41])  );
    wire logic pp_12_42;
    assign pp_12_42 = (select_e_12 & IN2[42] | select_2x_12 & IN2[41] | select_n2x_12 & (~ IN2[41]) | select_ne_12 & (~ IN2[42])  );
    wire logic pp_12_43;
    assign pp_12_43 = (select_e_12 & IN2[43] | select_2x_12 & IN2[42] | select_n2x_12 & (~ IN2[42]) | select_ne_12 & (~ IN2[43])  );
    wire logic pp_12_44;
    assign pp_12_44 = (select_e_12 & IN2[44] | select_2x_12 & IN2[43] | select_n2x_12 & (~ IN2[43]) | select_ne_12 & (~ IN2[44])  );
    wire logic pp_12_45;
    assign pp_12_45 = (select_e_12 & IN2[45] | select_2x_12 & IN2[44] | select_n2x_12 & (~ IN2[44]) | select_ne_12 & (~ IN2[45])  );
    wire logic pp_12_46;
    assign pp_12_46 = (select_e_12 & IN2[46] | select_2x_12 & IN2[45] | select_n2x_12 & (~ IN2[45]) | select_ne_12 & (~ IN2[46])  );
    wire logic pp_12_47;
    assign pp_12_47 = (select_e_12 & IN2[47] | select_2x_12 & IN2[46] | select_n2x_12 & (~ IN2[46]) | select_ne_12 & (~ IN2[47])  );
    wire logic pp_12_48;
    assign pp_12_48 = (select_e_12 & IN2[48] | select_2x_12 & IN2[47] | select_n2x_12 & (~ IN2[47]) | select_ne_12 & (~ IN2[48])  );
    wire logic pp_12_49;
    assign pp_12_49 = (select_e_12 & IN2[49] | select_2x_12 & IN2[48] | select_n2x_12 & (~ IN2[48]) | select_ne_12 & (~ IN2[49])  );
    wire logic pp_12_50;
    assign pp_12_50 = (select_e_12 & IN2[50] | select_2x_12 & IN2[49] | select_n2x_12 & (~ IN2[49]) | select_ne_12 & (~ IN2[50])  );
    wire logic pp_12_51;
    assign pp_12_51 = (select_e_12 & IN2[51] | select_2x_12 & IN2[50] | select_n2x_12 & (~ IN2[50]) | select_ne_12 & (~ IN2[51])  );
    wire logic pp_12_52;
    assign pp_12_52 = (select_e_12 & IN2[52] | select_2x_12 & IN2[51] | select_n2x_12 & (~ IN2[51]) | select_ne_12 & (~ IN2[52])  );
    wire logic pp_12_53;
    assign pp_12_53 = (select_e_12 & IN2[53] | select_2x_12 & IN2[52] | select_n2x_12 & (~ IN2[52]) | select_ne_12 & (~ IN2[53])  );
    wire logic pp_12_54;
    assign pp_12_54 = (select_e_12 & IN2[54] | select_2x_12 & IN2[53] | select_n2x_12 & (~ IN2[53]) | select_ne_12 & (~ IN2[54])  );
    wire logic pp_12_55;
    assign pp_12_55 = (select_e_12 & IN2[55] | select_2x_12 & IN2[54] | select_n2x_12 & (~ IN2[54]) | select_ne_12 & (~ IN2[55])  );
    wire logic pp_12_56;
    assign pp_12_56 = (select_e_12 & IN2[56] | select_2x_12 & IN2[55] | select_n2x_12 & (~ IN2[55]) | select_ne_12 & (~ IN2[56])  );
    wire logic pp_12_57;
    assign pp_12_57 = (select_e_12 & IN2[57] | select_2x_12 & IN2[56] | select_n2x_12 & (~ IN2[56]) | select_ne_12 & (~ IN2[57])  );
    wire logic pp_12_58;
    assign pp_12_58 = (select_e_12 & IN2[58] | select_2x_12 & IN2[57] | select_n2x_12 & (~ IN2[57]) | select_ne_12 & (~ IN2[58])  );
    wire logic pp_12_59;
    assign pp_12_59 = (select_e_12 & IN2[59] | select_2x_12 & IN2[58] | select_n2x_12 & (~ IN2[58]) | select_ne_12 & (~ IN2[59])  );
    wire logic pp_12_60;
    assign pp_12_60 = (select_e_12 & IN2[60] | select_2x_12 & IN2[59] | select_n2x_12 & (~ IN2[59]) | select_ne_12 & (~ IN2[60])  );
    wire logic pp_12_61;
    assign pp_12_61 = (select_e_12 & IN2[61] | select_2x_12 & IN2[60] | select_n2x_12 & (~ IN2[60]) | select_ne_12 & (~ IN2[61])  );
    wire logic pp_12_62;
    assign pp_12_62 = (select_e_12 & IN2[62] | select_2x_12 & IN2[61] | select_n2x_12 & (~ IN2[61]) | select_ne_12 & (~ IN2[62])  );
    wire logic pp_12_63;
    assign pp_12_63 = (select_e_12 & IN2[63] | select_2x_12 & IN2[62] | select_n2x_12 & (~ IN2[62]) | select_ne_12 & (~ IN2[63])  );
    wire logic pp_12_64;
    assign pp_12_64 = (select_e_12 & IN2[63] | select_2x_12 & IN2[63] | select_n2x_12 & (~ IN2[63]) | select_ne_12 & (~ IN2[63])  );
    wire logic pp_12_65;
    assign pp_12_65 = ~ (select_e_12 & IN2[63] | select_2x_12 & IN2[63] | select_n2x_12 & (~ IN2[63]) | select_ne_12 & (~ IN2[63])  );
    assign tcomp12 = select_ne_12 | select_n2x_12;
    
    // Signed Booth Radix-4 Partial Products Row 14
    wire logic select_e_13, select_ne_13, select_2x_13, tcomp13, select_n2x_13;
    assign select_e_13 = ((~ IN1[27]) & (IN1[26] ^ IN1[25]));
    assign select_ne_13 = IN1[27] &  (IN1[26] ^ IN1[25]);
    assign select_2x_13 = (~ IN1[27]) & IN1[26] & IN1[25];
    assign select_n2x_13 = IN1[27] & (~ IN1[26]) & (~ IN1[25]);
    wire logic pp_13_0;
    assign pp_13_0 = (select_e_13 & IN2[0] | select_2x_13 & 1'b0 | select_n2x_13 & 1'b1 | select_ne_13 & (~ IN2[0])  );
    wire logic pp_13_1;
    assign pp_13_1 = (select_e_13 & IN2[1] | select_2x_13 & IN2[0] | select_n2x_13 & (~ IN2[0]) | select_ne_13 & (~ IN2[1])  );
    wire logic pp_13_2;
    assign pp_13_2 = (select_e_13 & IN2[2] | select_2x_13 & IN2[1] | select_n2x_13 & (~ IN2[1]) | select_ne_13 & (~ IN2[2])  );
    wire logic pp_13_3;
    assign pp_13_3 = (select_e_13 & IN2[3] | select_2x_13 & IN2[2] | select_n2x_13 & (~ IN2[2]) | select_ne_13 & (~ IN2[3])  );
    wire logic pp_13_4;
    assign pp_13_4 = (select_e_13 & IN2[4] | select_2x_13 & IN2[3] | select_n2x_13 & (~ IN2[3]) | select_ne_13 & (~ IN2[4])  );
    wire logic pp_13_5;
    assign pp_13_5 = (select_e_13 & IN2[5] | select_2x_13 & IN2[4] | select_n2x_13 & (~ IN2[4]) | select_ne_13 & (~ IN2[5])  );
    wire logic pp_13_6;
    assign pp_13_6 = (select_e_13 & IN2[6] | select_2x_13 & IN2[5] | select_n2x_13 & (~ IN2[5]) | select_ne_13 & (~ IN2[6])  );
    wire logic pp_13_7;
    assign pp_13_7 = (select_e_13 & IN2[7] | select_2x_13 & IN2[6] | select_n2x_13 & (~ IN2[6]) | select_ne_13 & (~ IN2[7])  );
    wire logic pp_13_8;
    assign pp_13_8 = (select_e_13 & IN2[8] | select_2x_13 & IN2[7] | select_n2x_13 & (~ IN2[7]) | select_ne_13 & (~ IN2[8])  );
    wire logic pp_13_9;
    assign pp_13_9 = (select_e_13 & IN2[9] | select_2x_13 & IN2[8] | select_n2x_13 & (~ IN2[8]) | select_ne_13 & (~ IN2[9])  );
    wire logic pp_13_10;
    assign pp_13_10 = (select_e_13 & IN2[10] | select_2x_13 & IN2[9] | select_n2x_13 & (~ IN2[9]) | select_ne_13 & (~ IN2[10])  );
    wire logic pp_13_11;
    assign pp_13_11 = (select_e_13 & IN2[11] | select_2x_13 & IN2[10] | select_n2x_13 & (~ IN2[10]) | select_ne_13 & (~ IN2[11])  );
    wire logic pp_13_12;
    assign pp_13_12 = (select_e_13 & IN2[12] | select_2x_13 & IN2[11] | select_n2x_13 & (~ IN2[11]) | select_ne_13 & (~ IN2[12])  );
    wire logic pp_13_13;
    assign pp_13_13 = (select_e_13 & IN2[13] | select_2x_13 & IN2[12] | select_n2x_13 & (~ IN2[12]) | select_ne_13 & (~ IN2[13])  );
    wire logic pp_13_14;
    assign pp_13_14 = (select_e_13 & IN2[14] | select_2x_13 & IN2[13] | select_n2x_13 & (~ IN2[13]) | select_ne_13 & (~ IN2[14])  );
    wire logic pp_13_15;
    assign pp_13_15 = (select_e_13 & IN2[15] | select_2x_13 & IN2[14] | select_n2x_13 & (~ IN2[14]) | select_ne_13 & (~ IN2[15])  );
    wire logic pp_13_16;
    assign pp_13_16 = (select_e_13 & IN2[16] | select_2x_13 & IN2[15] | select_n2x_13 & (~ IN2[15]) | select_ne_13 & (~ IN2[16])  );
    wire logic pp_13_17;
    assign pp_13_17 = (select_e_13 & IN2[17] | select_2x_13 & IN2[16] | select_n2x_13 & (~ IN2[16]) | select_ne_13 & (~ IN2[17])  );
    wire logic pp_13_18;
    assign pp_13_18 = (select_e_13 & IN2[18] | select_2x_13 & IN2[17] | select_n2x_13 & (~ IN2[17]) | select_ne_13 & (~ IN2[18])  );
    wire logic pp_13_19;
    assign pp_13_19 = (select_e_13 & IN2[19] | select_2x_13 & IN2[18] | select_n2x_13 & (~ IN2[18]) | select_ne_13 & (~ IN2[19])  );
    wire logic pp_13_20;
    assign pp_13_20 = (select_e_13 & IN2[20] | select_2x_13 & IN2[19] | select_n2x_13 & (~ IN2[19]) | select_ne_13 & (~ IN2[20])  );
    wire logic pp_13_21;
    assign pp_13_21 = (select_e_13 & IN2[21] | select_2x_13 & IN2[20] | select_n2x_13 & (~ IN2[20]) | select_ne_13 & (~ IN2[21])  );
    wire logic pp_13_22;
    assign pp_13_22 = (select_e_13 & IN2[22] | select_2x_13 & IN2[21] | select_n2x_13 & (~ IN2[21]) | select_ne_13 & (~ IN2[22])  );
    wire logic pp_13_23;
    assign pp_13_23 = (select_e_13 & IN2[23] | select_2x_13 & IN2[22] | select_n2x_13 & (~ IN2[22]) | select_ne_13 & (~ IN2[23])  );
    wire logic pp_13_24;
    assign pp_13_24 = (select_e_13 & IN2[24] | select_2x_13 & IN2[23] | select_n2x_13 & (~ IN2[23]) | select_ne_13 & (~ IN2[24])  );
    wire logic pp_13_25;
    assign pp_13_25 = (select_e_13 & IN2[25] | select_2x_13 & IN2[24] | select_n2x_13 & (~ IN2[24]) | select_ne_13 & (~ IN2[25])  );
    wire logic pp_13_26;
    assign pp_13_26 = (select_e_13 & IN2[26] | select_2x_13 & IN2[25] | select_n2x_13 & (~ IN2[25]) | select_ne_13 & (~ IN2[26])  );
    wire logic pp_13_27;
    assign pp_13_27 = (select_e_13 & IN2[27] | select_2x_13 & IN2[26] | select_n2x_13 & (~ IN2[26]) | select_ne_13 & (~ IN2[27])  );
    wire logic pp_13_28;
    assign pp_13_28 = (select_e_13 & IN2[28] | select_2x_13 & IN2[27] | select_n2x_13 & (~ IN2[27]) | select_ne_13 & (~ IN2[28])  );
    wire logic pp_13_29;
    assign pp_13_29 = (select_e_13 & IN2[29] | select_2x_13 & IN2[28] | select_n2x_13 & (~ IN2[28]) | select_ne_13 & (~ IN2[29])  );
    wire logic pp_13_30;
    assign pp_13_30 = (select_e_13 & IN2[30] | select_2x_13 & IN2[29] | select_n2x_13 & (~ IN2[29]) | select_ne_13 & (~ IN2[30])  );
    wire logic pp_13_31;
    assign pp_13_31 = (select_e_13 & IN2[31] | select_2x_13 & IN2[30] | select_n2x_13 & (~ IN2[30]) | select_ne_13 & (~ IN2[31])  );
    wire logic pp_13_32;
    assign pp_13_32 = (select_e_13 & IN2[32] | select_2x_13 & IN2[31] | select_n2x_13 & (~ IN2[31]) | select_ne_13 & (~ IN2[32])  );
    wire logic pp_13_33;
    assign pp_13_33 = (select_e_13 & IN2[33] | select_2x_13 & IN2[32] | select_n2x_13 & (~ IN2[32]) | select_ne_13 & (~ IN2[33])  );
    wire logic pp_13_34;
    assign pp_13_34 = (select_e_13 & IN2[34] | select_2x_13 & IN2[33] | select_n2x_13 & (~ IN2[33]) | select_ne_13 & (~ IN2[34])  );
    wire logic pp_13_35;
    assign pp_13_35 = (select_e_13 & IN2[35] | select_2x_13 & IN2[34] | select_n2x_13 & (~ IN2[34]) | select_ne_13 & (~ IN2[35])  );
    wire logic pp_13_36;
    assign pp_13_36 = (select_e_13 & IN2[36] | select_2x_13 & IN2[35] | select_n2x_13 & (~ IN2[35]) | select_ne_13 & (~ IN2[36])  );
    wire logic pp_13_37;
    assign pp_13_37 = (select_e_13 & IN2[37] | select_2x_13 & IN2[36] | select_n2x_13 & (~ IN2[36]) | select_ne_13 & (~ IN2[37])  );
    wire logic pp_13_38;
    assign pp_13_38 = (select_e_13 & IN2[38] | select_2x_13 & IN2[37] | select_n2x_13 & (~ IN2[37]) | select_ne_13 & (~ IN2[38])  );
    wire logic pp_13_39;
    assign pp_13_39 = (select_e_13 & IN2[39] | select_2x_13 & IN2[38] | select_n2x_13 & (~ IN2[38]) | select_ne_13 & (~ IN2[39])  );
    wire logic pp_13_40;
    assign pp_13_40 = (select_e_13 & IN2[40] | select_2x_13 & IN2[39] | select_n2x_13 & (~ IN2[39]) | select_ne_13 & (~ IN2[40])  );
    wire logic pp_13_41;
    assign pp_13_41 = (select_e_13 & IN2[41] | select_2x_13 & IN2[40] | select_n2x_13 & (~ IN2[40]) | select_ne_13 & (~ IN2[41])  );
    wire logic pp_13_42;
    assign pp_13_42 = (select_e_13 & IN2[42] | select_2x_13 & IN2[41] | select_n2x_13 & (~ IN2[41]) | select_ne_13 & (~ IN2[42])  );
    wire logic pp_13_43;
    assign pp_13_43 = (select_e_13 & IN2[43] | select_2x_13 & IN2[42] | select_n2x_13 & (~ IN2[42]) | select_ne_13 & (~ IN2[43])  );
    wire logic pp_13_44;
    assign pp_13_44 = (select_e_13 & IN2[44] | select_2x_13 & IN2[43] | select_n2x_13 & (~ IN2[43]) | select_ne_13 & (~ IN2[44])  );
    wire logic pp_13_45;
    assign pp_13_45 = (select_e_13 & IN2[45] | select_2x_13 & IN2[44] | select_n2x_13 & (~ IN2[44]) | select_ne_13 & (~ IN2[45])  );
    wire logic pp_13_46;
    assign pp_13_46 = (select_e_13 & IN2[46] | select_2x_13 & IN2[45] | select_n2x_13 & (~ IN2[45]) | select_ne_13 & (~ IN2[46])  );
    wire logic pp_13_47;
    assign pp_13_47 = (select_e_13 & IN2[47] | select_2x_13 & IN2[46] | select_n2x_13 & (~ IN2[46]) | select_ne_13 & (~ IN2[47])  );
    wire logic pp_13_48;
    assign pp_13_48 = (select_e_13 & IN2[48] | select_2x_13 & IN2[47] | select_n2x_13 & (~ IN2[47]) | select_ne_13 & (~ IN2[48])  );
    wire logic pp_13_49;
    assign pp_13_49 = (select_e_13 & IN2[49] | select_2x_13 & IN2[48] | select_n2x_13 & (~ IN2[48]) | select_ne_13 & (~ IN2[49])  );
    wire logic pp_13_50;
    assign pp_13_50 = (select_e_13 & IN2[50] | select_2x_13 & IN2[49] | select_n2x_13 & (~ IN2[49]) | select_ne_13 & (~ IN2[50])  );
    wire logic pp_13_51;
    assign pp_13_51 = (select_e_13 & IN2[51] | select_2x_13 & IN2[50] | select_n2x_13 & (~ IN2[50]) | select_ne_13 & (~ IN2[51])  );
    wire logic pp_13_52;
    assign pp_13_52 = (select_e_13 & IN2[52] | select_2x_13 & IN2[51] | select_n2x_13 & (~ IN2[51]) | select_ne_13 & (~ IN2[52])  );
    wire logic pp_13_53;
    assign pp_13_53 = (select_e_13 & IN2[53] | select_2x_13 & IN2[52] | select_n2x_13 & (~ IN2[52]) | select_ne_13 & (~ IN2[53])  );
    wire logic pp_13_54;
    assign pp_13_54 = (select_e_13 & IN2[54] | select_2x_13 & IN2[53] | select_n2x_13 & (~ IN2[53]) | select_ne_13 & (~ IN2[54])  );
    wire logic pp_13_55;
    assign pp_13_55 = (select_e_13 & IN2[55] | select_2x_13 & IN2[54] | select_n2x_13 & (~ IN2[54]) | select_ne_13 & (~ IN2[55])  );
    wire logic pp_13_56;
    assign pp_13_56 = (select_e_13 & IN2[56] | select_2x_13 & IN2[55] | select_n2x_13 & (~ IN2[55]) | select_ne_13 & (~ IN2[56])  );
    wire logic pp_13_57;
    assign pp_13_57 = (select_e_13 & IN2[57] | select_2x_13 & IN2[56] | select_n2x_13 & (~ IN2[56]) | select_ne_13 & (~ IN2[57])  );
    wire logic pp_13_58;
    assign pp_13_58 = (select_e_13 & IN2[58] | select_2x_13 & IN2[57] | select_n2x_13 & (~ IN2[57]) | select_ne_13 & (~ IN2[58])  );
    wire logic pp_13_59;
    assign pp_13_59 = (select_e_13 & IN2[59] | select_2x_13 & IN2[58] | select_n2x_13 & (~ IN2[58]) | select_ne_13 & (~ IN2[59])  );
    wire logic pp_13_60;
    assign pp_13_60 = (select_e_13 & IN2[60] | select_2x_13 & IN2[59] | select_n2x_13 & (~ IN2[59]) | select_ne_13 & (~ IN2[60])  );
    wire logic pp_13_61;
    assign pp_13_61 = (select_e_13 & IN2[61] | select_2x_13 & IN2[60] | select_n2x_13 & (~ IN2[60]) | select_ne_13 & (~ IN2[61])  );
    wire logic pp_13_62;
    assign pp_13_62 = (select_e_13 & IN2[62] | select_2x_13 & IN2[61] | select_n2x_13 & (~ IN2[61]) | select_ne_13 & (~ IN2[62])  );
    wire logic pp_13_63;
    assign pp_13_63 = (select_e_13 & IN2[63] | select_2x_13 & IN2[62] | select_n2x_13 & (~ IN2[62]) | select_ne_13 & (~ IN2[63])  );
    wire logic pp_13_64;
    assign pp_13_64 = (select_e_13 & IN2[63] | select_2x_13 & IN2[63] | select_n2x_13 & (~ IN2[63]) | select_ne_13 & (~ IN2[63])  );
    wire logic pp_13_65;
    assign pp_13_65 = ~ (select_e_13 & IN2[63] | select_2x_13 & IN2[63] | select_n2x_13 & (~ IN2[63]) | select_ne_13 & (~ IN2[63])  );
    assign tcomp13 = select_ne_13 | select_n2x_13;
    
    // Signed Booth Radix-4 Partial Products Row 15
    wire logic select_e_14, select_ne_14, select_2x_14, tcomp14, select_n2x_14;
    assign select_e_14 = ((~ IN1[29]) & (IN1[28] ^ IN1[27]));
    assign select_ne_14 = IN1[29] &  (IN1[28] ^ IN1[27]);
    assign select_2x_14 = (~ IN1[29]) & IN1[28] & IN1[27];
    assign select_n2x_14 = IN1[29] & (~ IN1[28]) & (~ IN1[27]);
    wire logic pp_14_0;
    assign pp_14_0 = (select_e_14 & IN2[0] | select_2x_14 & 1'b0 | select_n2x_14 & 1'b1 | select_ne_14 & (~ IN2[0])  );
    wire logic pp_14_1;
    assign pp_14_1 = (select_e_14 & IN2[1] | select_2x_14 & IN2[0] | select_n2x_14 & (~ IN2[0]) | select_ne_14 & (~ IN2[1])  );
    wire logic pp_14_2;
    assign pp_14_2 = (select_e_14 & IN2[2] | select_2x_14 & IN2[1] | select_n2x_14 & (~ IN2[1]) | select_ne_14 & (~ IN2[2])  );
    wire logic pp_14_3;
    assign pp_14_3 = (select_e_14 & IN2[3] | select_2x_14 & IN2[2] | select_n2x_14 & (~ IN2[2]) | select_ne_14 & (~ IN2[3])  );
    wire logic pp_14_4;
    assign pp_14_4 = (select_e_14 & IN2[4] | select_2x_14 & IN2[3] | select_n2x_14 & (~ IN2[3]) | select_ne_14 & (~ IN2[4])  );
    wire logic pp_14_5;
    assign pp_14_5 = (select_e_14 & IN2[5] | select_2x_14 & IN2[4] | select_n2x_14 & (~ IN2[4]) | select_ne_14 & (~ IN2[5])  );
    wire logic pp_14_6;
    assign pp_14_6 = (select_e_14 & IN2[6] | select_2x_14 & IN2[5] | select_n2x_14 & (~ IN2[5]) | select_ne_14 & (~ IN2[6])  );
    wire logic pp_14_7;
    assign pp_14_7 = (select_e_14 & IN2[7] | select_2x_14 & IN2[6] | select_n2x_14 & (~ IN2[6]) | select_ne_14 & (~ IN2[7])  );
    wire logic pp_14_8;
    assign pp_14_8 = (select_e_14 & IN2[8] | select_2x_14 & IN2[7] | select_n2x_14 & (~ IN2[7]) | select_ne_14 & (~ IN2[8])  );
    wire logic pp_14_9;
    assign pp_14_9 = (select_e_14 & IN2[9] | select_2x_14 & IN2[8] | select_n2x_14 & (~ IN2[8]) | select_ne_14 & (~ IN2[9])  );
    wire logic pp_14_10;
    assign pp_14_10 = (select_e_14 & IN2[10] | select_2x_14 & IN2[9] | select_n2x_14 & (~ IN2[9]) | select_ne_14 & (~ IN2[10])  );
    wire logic pp_14_11;
    assign pp_14_11 = (select_e_14 & IN2[11] | select_2x_14 & IN2[10] | select_n2x_14 & (~ IN2[10]) | select_ne_14 & (~ IN2[11])  );
    wire logic pp_14_12;
    assign pp_14_12 = (select_e_14 & IN2[12] | select_2x_14 & IN2[11] | select_n2x_14 & (~ IN2[11]) | select_ne_14 & (~ IN2[12])  );
    wire logic pp_14_13;
    assign pp_14_13 = (select_e_14 & IN2[13] | select_2x_14 & IN2[12] | select_n2x_14 & (~ IN2[12]) | select_ne_14 & (~ IN2[13])  );
    wire logic pp_14_14;
    assign pp_14_14 = (select_e_14 & IN2[14] | select_2x_14 & IN2[13] | select_n2x_14 & (~ IN2[13]) | select_ne_14 & (~ IN2[14])  );
    wire logic pp_14_15;
    assign pp_14_15 = (select_e_14 & IN2[15] | select_2x_14 & IN2[14] | select_n2x_14 & (~ IN2[14]) | select_ne_14 & (~ IN2[15])  );
    wire logic pp_14_16;
    assign pp_14_16 = (select_e_14 & IN2[16] | select_2x_14 & IN2[15] | select_n2x_14 & (~ IN2[15]) | select_ne_14 & (~ IN2[16])  );
    wire logic pp_14_17;
    assign pp_14_17 = (select_e_14 & IN2[17] | select_2x_14 & IN2[16] | select_n2x_14 & (~ IN2[16]) | select_ne_14 & (~ IN2[17])  );
    wire logic pp_14_18;
    assign pp_14_18 = (select_e_14 & IN2[18] | select_2x_14 & IN2[17] | select_n2x_14 & (~ IN2[17]) | select_ne_14 & (~ IN2[18])  );
    wire logic pp_14_19;
    assign pp_14_19 = (select_e_14 & IN2[19] | select_2x_14 & IN2[18] | select_n2x_14 & (~ IN2[18]) | select_ne_14 & (~ IN2[19])  );
    wire logic pp_14_20;
    assign pp_14_20 = (select_e_14 & IN2[20] | select_2x_14 & IN2[19] | select_n2x_14 & (~ IN2[19]) | select_ne_14 & (~ IN2[20])  );
    wire logic pp_14_21;
    assign pp_14_21 = (select_e_14 & IN2[21] | select_2x_14 & IN2[20] | select_n2x_14 & (~ IN2[20]) | select_ne_14 & (~ IN2[21])  );
    wire logic pp_14_22;
    assign pp_14_22 = (select_e_14 & IN2[22] | select_2x_14 & IN2[21] | select_n2x_14 & (~ IN2[21]) | select_ne_14 & (~ IN2[22])  );
    wire logic pp_14_23;
    assign pp_14_23 = (select_e_14 & IN2[23] | select_2x_14 & IN2[22] | select_n2x_14 & (~ IN2[22]) | select_ne_14 & (~ IN2[23])  );
    wire logic pp_14_24;
    assign pp_14_24 = (select_e_14 & IN2[24] | select_2x_14 & IN2[23] | select_n2x_14 & (~ IN2[23]) | select_ne_14 & (~ IN2[24])  );
    wire logic pp_14_25;
    assign pp_14_25 = (select_e_14 & IN2[25] | select_2x_14 & IN2[24] | select_n2x_14 & (~ IN2[24]) | select_ne_14 & (~ IN2[25])  );
    wire logic pp_14_26;
    assign pp_14_26 = (select_e_14 & IN2[26] | select_2x_14 & IN2[25] | select_n2x_14 & (~ IN2[25]) | select_ne_14 & (~ IN2[26])  );
    wire logic pp_14_27;
    assign pp_14_27 = (select_e_14 & IN2[27] | select_2x_14 & IN2[26] | select_n2x_14 & (~ IN2[26]) | select_ne_14 & (~ IN2[27])  );
    wire logic pp_14_28;
    assign pp_14_28 = (select_e_14 & IN2[28] | select_2x_14 & IN2[27] | select_n2x_14 & (~ IN2[27]) | select_ne_14 & (~ IN2[28])  );
    wire logic pp_14_29;
    assign pp_14_29 = (select_e_14 & IN2[29] | select_2x_14 & IN2[28] | select_n2x_14 & (~ IN2[28]) | select_ne_14 & (~ IN2[29])  );
    wire logic pp_14_30;
    assign pp_14_30 = (select_e_14 & IN2[30] | select_2x_14 & IN2[29] | select_n2x_14 & (~ IN2[29]) | select_ne_14 & (~ IN2[30])  );
    wire logic pp_14_31;
    assign pp_14_31 = (select_e_14 & IN2[31] | select_2x_14 & IN2[30] | select_n2x_14 & (~ IN2[30]) | select_ne_14 & (~ IN2[31])  );
    wire logic pp_14_32;
    assign pp_14_32 = (select_e_14 & IN2[32] | select_2x_14 & IN2[31] | select_n2x_14 & (~ IN2[31]) | select_ne_14 & (~ IN2[32])  );
    wire logic pp_14_33;
    assign pp_14_33 = (select_e_14 & IN2[33] | select_2x_14 & IN2[32] | select_n2x_14 & (~ IN2[32]) | select_ne_14 & (~ IN2[33])  );
    wire logic pp_14_34;
    assign pp_14_34 = (select_e_14 & IN2[34] | select_2x_14 & IN2[33] | select_n2x_14 & (~ IN2[33]) | select_ne_14 & (~ IN2[34])  );
    wire logic pp_14_35;
    assign pp_14_35 = (select_e_14 & IN2[35] | select_2x_14 & IN2[34] | select_n2x_14 & (~ IN2[34]) | select_ne_14 & (~ IN2[35])  );
    wire logic pp_14_36;
    assign pp_14_36 = (select_e_14 & IN2[36] | select_2x_14 & IN2[35] | select_n2x_14 & (~ IN2[35]) | select_ne_14 & (~ IN2[36])  );
    wire logic pp_14_37;
    assign pp_14_37 = (select_e_14 & IN2[37] | select_2x_14 & IN2[36] | select_n2x_14 & (~ IN2[36]) | select_ne_14 & (~ IN2[37])  );
    wire logic pp_14_38;
    assign pp_14_38 = (select_e_14 & IN2[38] | select_2x_14 & IN2[37] | select_n2x_14 & (~ IN2[37]) | select_ne_14 & (~ IN2[38])  );
    wire logic pp_14_39;
    assign pp_14_39 = (select_e_14 & IN2[39] | select_2x_14 & IN2[38] | select_n2x_14 & (~ IN2[38]) | select_ne_14 & (~ IN2[39])  );
    wire logic pp_14_40;
    assign pp_14_40 = (select_e_14 & IN2[40] | select_2x_14 & IN2[39] | select_n2x_14 & (~ IN2[39]) | select_ne_14 & (~ IN2[40])  );
    wire logic pp_14_41;
    assign pp_14_41 = (select_e_14 & IN2[41] | select_2x_14 & IN2[40] | select_n2x_14 & (~ IN2[40]) | select_ne_14 & (~ IN2[41])  );
    wire logic pp_14_42;
    assign pp_14_42 = (select_e_14 & IN2[42] | select_2x_14 & IN2[41] | select_n2x_14 & (~ IN2[41]) | select_ne_14 & (~ IN2[42])  );
    wire logic pp_14_43;
    assign pp_14_43 = (select_e_14 & IN2[43] | select_2x_14 & IN2[42] | select_n2x_14 & (~ IN2[42]) | select_ne_14 & (~ IN2[43])  );
    wire logic pp_14_44;
    assign pp_14_44 = (select_e_14 & IN2[44] | select_2x_14 & IN2[43] | select_n2x_14 & (~ IN2[43]) | select_ne_14 & (~ IN2[44])  );
    wire logic pp_14_45;
    assign pp_14_45 = (select_e_14 & IN2[45] | select_2x_14 & IN2[44] | select_n2x_14 & (~ IN2[44]) | select_ne_14 & (~ IN2[45])  );
    wire logic pp_14_46;
    assign pp_14_46 = (select_e_14 & IN2[46] | select_2x_14 & IN2[45] | select_n2x_14 & (~ IN2[45]) | select_ne_14 & (~ IN2[46])  );
    wire logic pp_14_47;
    assign pp_14_47 = (select_e_14 & IN2[47] | select_2x_14 & IN2[46] | select_n2x_14 & (~ IN2[46]) | select_ne_14 & (~ IN2[47])  );
    wire logic pp_14_48;
    assign pp_14_48 = (select_e_14 & IN2[48] | select_2x_14 & IN2[47] | select_n2x_14 & (~ IN2[47]) | select_ne_14 & (~ IN2[48])  );
    wire logic pp_14_49;
    assign pp_14_49 = (select_e_14 & IN2[49] | select_2x_14 & IN2[48] | select_n2x_14 & (~ IN2[48]) | select_ne_14 & (~ IN2[49])  );
    wire logic pp_14_50;
    assign pp_14_50 = (select_e_14 & IN2[50] | select_2x_14 & IN2[49] | select_n2x_14 & (~ IN2[49]) | select_ne_14 & (~ IN2[50])  );
    wire logic pp_14_51;
    assign pp_14_51 = (select_e_14 & IN2[51] | select_2x_14 & IN2[50] | select_n2x_14 & (~ IN2[50]) | select_ne_14 & (~ IN2[51])  );
    wire logic pp_14_52;
    assign pp_14_52 = (select_e_14 & IN2[52] | select_2x_14 & IN2[51] | select_n2x_14 & (~ IN2[51]) | select_ne_14 & (~ IN2[52])  );
    wire logic pp_14_53;
    assign pp_14_53 = (select_e_14 & IN2[53] | select_2x_14 & IN2[52] | select_n2x_14 & (~ IN2[52]) | select_ne_14 & (~ IN2[53])  );
    wire logic pp_14_54;
    assign pp_14_54 = (select_e_14 & IN2[54] | select_2x_14 & IN2[53] | select_n2x_14 & (~ IN2[53]) | select_ne_14 & (~ IN2[54])  );
    wire logic pp_14_55;
    assign pp_14_55 = (select_e_14 & IN2[55] | select_2x_14 & IN2[54] | select_n2x_14 & (~ IN2[54]) | select_ne_14 & (~ IN2[55])  );
    wire logic pp_14_56;
    assign pp_14_56 = (select_e_14 & IN2[56] | select_2x_14 & IN2[55] | select_n2x_14 & (~ IN2[55]) | select_ne_14 & (~ IN2[56])  );
    wire logic pp_14_57;
    assign pp_14_57 = (select_e_14 & IN2[57] | select_2x_14 & IN2[56] | select_n2x_14 & (~ IN2[56]) | select_ne_14 & (~ IN2[57])  );
    wire logic pp_14_58;
    assign pp_14_58 = (select_e_14 & IN2[58] | select_2x_14 & IN2[57] | select_n2x_14 & (~ IN2[57]) | select_ne_14 & (~ IN2[58])  );
    wire logic pp_14_59;
    assign pp_14_59 = (select_e_14 & IN2[59] | select_2x_14 & IN2[58] | select_n2x_14 & (~ IN2[58]) | select_ne_14 & (~ IN2[59])  );
    wire logic pp_14_60;
    assign pp_14_60 = (select_e_14 & IN2[60] | select_2x_14 & IN2[59] | select_n2x_14 & (~ IN2[59]) | select_ne_14 & (~ IN2[60])  );
    wire logic pp_14_61;
    assign pp_14_61 = (select_e_14 & IN2[61] | select_2x_14 & IN2[60] | select_n2x_14 & (~ IN2[60]) | select_ne_14 & (~ IN2[61])  );
    wire logic pp_14_62;
    assign pp_14_62 = (select_e_14 & IN2[62] | select_2x_14 & IN2[61] | select_n2x_14 & (~ IN2[61]) | select_ne_14 & (~ IN2[62])  );
    wire logic pp_14_63;
    assign pp_14_63 = (select_e_14 & IN2[63] | select_2x_14 & IN2[62] | select_n2x_14 & (~ IN2[62]) | select_ne_14 & (~ IN2[63])  );
    wire logic pp_14_64;
    assign pp_14_64 = (select_e_14 & IN2[63] | select_2x_14 & IN2[63] | select_n2x_14 & (~ IN2[63]) | select_ne_14 & (~ IN2[63])  );
    wire logic pp_14_65;
    assign pp_14_65 = ~ (select_e_14 & IN2[63] | select_2x_14 & IN2[63] | select_n2x_14 & (~ IN2[63]) | select_ne_14 & (~ IN2[63])  );
    assign tcomp14 = select_ne_14 | select_n2x_14;
    
    // Signed Booth Radix-4 Partial Products Row 16
    wire logic select_e_15, select_ne_15, select_2x_15, tcomp15, select_n2x_15;
    assign select_e_15 = ((~ IN1[31]) & (IN1[30] ^ IN1[29]));
    assign select_ne_15 = IN1[31] &  (IN1[30] ^ IN1[29]);
    assign select_2x_15 = (~ IN1[31]) & IN1[30] & IN1[29];
    assign select_n2x_15 = IN1[31] & (~ IN1[30]) & (~ IN1[29]);
    wire logic pp_15_0;
    assign pp_15_0 = (select_e_15 & IN2[0] | select_2x_15 & 1'b0 | select_n2x_15 & 1'b1 | select_ne_15 & (~ IN2[0])  );
    wire logic pp_15_1;
    assign pp_15_1 = (select_e_15 & IN2[1] | select_2x_15 & IN2[0] | select_n2x_15 & (~ IN2[0]) | select_ne_15 & (~ IN2[1])  );
    wire logic pp_15_2;
    assign pp_15_2 = (select_e_15 & IN2[2] | select_2x_15 & IN2[1] | select_n2x_15 & (~ IN2[1]) | select_ne_15 & (~ IN2[2])  );
    wire logic pp_15_3;
    assign pp_15_3 = (select_e_15 & IN2[3] | select_2x_15 & IN2[2] | select_n2x_15 & (~ IN2[2]) | select_ne_15 & (~ IN2[3])  );
    wire logic pp_15_4;
    assign pp_15_4 = (select_e_15 & IN2[4] | select_2x_15 & IN2[3] | select_n2x_15 & (~ IN2[3]) | select_ne_15 & (~ IN2[4])  );
    wire logic pp_15_5;
    assign pp_15_5 = (select_e_15 & IN2[5] | select_2x_15 & IN2[4] | select_n2x_15 & (~ IN2[4]) | select_ne_15 & (~ IN2[5])  );
    wire logic pp_15_6;
    assign pp_15_6 = (select_e_15 & IN2[6] | select_2x_15 & IN2[5] | select_n2x_15 & (~ IN2[5]) | select_ne_15 & (~ IN2[6])  );
    wire logic pp_15_7;
    assign pp_15_7 = (select_e_15 & IN2[7] | select_2x_15 & IN2[6] | select_n2x_15 & (~ IN2[6]) | select_ne_15 & (~ IN2[7])  );
    wire logic pp_15_8;
    assign pp_15_8 = (select_e_15 & IN2[8] | select_2x_15 & IN2[7] | select_n2x_15 & (~ IN2[7]) | select_ne_15 & (~ IN2[8])  );
    wire logic pp_15_9;
    assign pp_15_9 = (select_e_15 & IN2[9] | select_2x_15 & IN2[8] | select_n2x_15 & (~ IN2[8]) | select_ne_15 & (~ IN2[9])  );
    wire logic pp_15_10;
    assign pp_15_10 = (select_e_15 & IN2[10] | select_2x_15 & IN2[9] | select_n2x_15 & (~ IN2[9]) | select_ne_15 & (~ IN2[10])  );
    wire logic pp_15_11;
    assign pp_15_11 = (select_e_15 & IN2[11] | select_2x_15 & IN2[10] | select_n2x_15 & (~ IN2[10]) | select_ne_15 & (~ IN2[11])  );
    wire logic pp_15_12;
    assign pp_15_12 = (select_e_15 & IN2[12] | select_2x_15 & IN2[11] | select_n2x_15 & (~ IN2[11]) | select_ne_15 & (~ IN2[12])  );
    wire logic pp_15_13;
    assign pp_15_13 = (select_e_15 & IN2[13] | select_2x_15 & IN2[12] | select_n2x_15 & (~ IN2[12]) | select_ne_15 & (~ IN2[13])  );
    wire logic pp_15_14;
    assign pp_15_14 = (select_e_15 & IN2[14] | select_2x_15 & IN2[13] | select_n2x_15 & (~ IN2[13]) | select_ne_15 & (~ IN2[14])  );
    wire logic pp_15_15;
    assign pp_15_15 = (select_e_15 & IN2[15] | select_2x_15 & IN2[14] | select_n2x_15 & (~ IN2[14]) | select_ne_15 & (~ IN2[15])  );
    wire logic pp_15_16;
    assign pp_15_16 = (select_e_15 & IN2[16] | select_2x_15 & IN2[15] | select_n2x_15 & (~ IN2[15]) | select_ne_15 & (~ IN2[16])  );
    wire logic pp_15_17;
    assign pp_15_17 = (select_e_15 & IN2[17] | select_2x_15 & IN2[16] | select_n2x_15 & (~ IN2[16]) | select_ne_15 & (~ IN2[17])  );
    wire logic pp_15_18;
    assign pp_15_18 = (select_e_15 & IN2[18] | select_2x_15 & IN2[17] | select_n2x_15 & (~ IN2[17]) | select_ne_15 & (~ IN2[18])  );
    wire logic pp_15_19;
    assign pp_15_19 = (select_e_15 & IN2[19] | select_2x_15 & IN2[18] | select_n2x_15 & (~ IN2[18]) | select_ne_15 & (~ IN2[19])  );
    wire logic pp_15_20;
    assign pp_15_20 = (select_e_15 & IN2[20] | select_2x_15 & IN2[19] | select_n2x_15 & (~ IN2[19]) | select_ne_15 & (~ IN2[20])  );
    wire logic pp_15_21;
    assign pp_15_21 = (select_e_15 & IN2[21] | select_2x_15 & IN2[20] | select_n2x_15 & (~ IN2[20]) | select_ne_15 & (~ IN2[21])  );
    wire logic pp_15_22;
    assign pp_15_22 = (select_e_15 & IN2[22] | select_2x_15 & IN2[21] | select_n2x_15 & (~ IN2[21]) | select_ne_15 & (~ IN2[22])  );
    wire logic pp_15_23;
    assign pp_15_23 = (select_e_15 & IN2[23] | select_2x_15 & IN2[22] | select_n2x_15 & (~ IN2[22]) | select_ne_15 & (~ IN2[23])  );
    wire logic pp_15_24;
    assign pp_15_24 = (select_e_15 & IN2[24] | select_2x_15 & IN2[23] | select_n2x_15 & (~ IN2[23]) | select_ne_15 & (~ IN2[24])  );
    wire logic pp_15_25;
    assign pp_15_25 = (select_e_15 & IN2[25] | select_2x_15 & IN2[24] | select_n2x_15 & (~ IN2[24]) | select_ne_15 & (~ IN2[25])  );
    wire logic pp_15_26;
    assign pp_15_26 = (select_e_15 & IN2[26] | select_2x_15 & IN2[25] | select_n2x_15 & (~ IN2[25]) | select_ne_15 & (~ IN2[26])  );
    wire logic pp_15_27;
    assign pp_15_27 = (select_e_15 & IN2[27] | select_2x_15 & IN2[26] | select_n2x_15 & (~ IN2[26]) | select_ne_15 & (~ IN2[27])  );
    wire logic pp_15_28;
    assign pp_15_28 = (select_e_15 & IN2[28] | select_2x_15 & IN2[27] | select_n2x_15 & (~ IN2[27]) | select_ne_15 & (~ IN2[28])  );
    wire logic pp_15_29;
    assign pp_15_29 = (select_e_15 & IN2[29] | select_2x_15 & IN2[28] | select_n2x_15 & (~ IN2[28]) | select_ne_15 & (~ IN2[29])  );
    wire logic pp_15_30;
    assign pp_15_30 = (select_e_15 & IN2[30] | select_2x_15 & IN2[29] | select_n2x_15 & (~ IN2[29]) | select_ne_15 & (~ IN2[30])  );
    wire logic pp_15_31;
    assign pp_15_31 = (select_e_15 & IN2[31] | select_2x_15 & IN2[30] | select_n2x_15 & (~ IN2[30]) | select_ne_15 & (~ IN2[31])  );
    wire logic pp_15_32;
    assign pp_15_32 = (select_e_15 & IN2[32] | select_2x_15 & IN2[31] | select_n2x_15 & (~ IN2[31]) | select_ne_15 & (~ IN2[32])  );
    wire logic pp_15_33;
    assign pp_15_33 = (select_e_15 & IN2[33] | select_2x_15 & IN2[32] | select_n2x_15 & (~ IN2[32]) | select_ne_15 & (~ IN2[33])  );
    wire logic pp_15_34;
    assign pp_15_34 = (select_e_15 & IN2[34] | select_2x_15 & IN2[33] | select_n2x_15 & (~ IN2[33]) | select_ne_15 & (~ IN2[34])  );
    wire logic pp_15_35;
    assign pp_15_35 = (select_e_15 & IN2[35] | select_2x_15 & IN2[34] | select_n2x_15 & (~ IN2[34]) | select_ne_15 & (~ IN2[35])  );
    wire logic pp_15_36;
    assign pp_15_36 = (select_e_15 & IN2[36] | select_2x_15 & IN2[35] | select_n2x_15 & (~ IN2[35]) | select_ne_15 & (~ IN2[36])  );
    wire logic pp_15_37;
    assign pp_15_37 = (select_e_15 & IN2[37] | select_2x_15 & IN2[36] | select_n2x_15 & (~ IN2[36]) | select_ne_15 & (~ IN2[37])  );
    wire logic pp_15_38;
    assign pp_15_38 = (select_e_15 & IN2[38] | select_2x_15 & IN2[37] | select_n2x_15 & (~ IN2[37]) | select_ne_15 & (~ IN2[38])  );
    wire logic pp_15_39;
    assign pp_15_39 = (select_e_15 & IN2[39] | select_2x_15 & IN2[38] | select_n2x_15 & (~ IN2[38]) | select_ne_15 & (~ IN2[39])  );
    wire logic pp_15_40;
    assign pp_15_40 = (select_e_15 & IN2[40] | select_2x_15 & IN2[39] | select_n2x_15 & (~ IN2[39]) | select_ne_15 & (~ IN2[40])  );
    wire logic pp_15_41;
    assign pp_15_41 = (select_e_15 & IN2[41] | select_2x_15 & IN2[40] | select_n2x_15 & (~ IN2[40]) | select_ne_15 & (~ IN2[41])  );
    wire logic pp_15_42;
    assign pp_15_42 = (select_e_15 & IN2[42] | select_2x_15 & IN2[41] | select_n2x_15 & (~ IN2[41]) | select_ne_15 & (~ IN2[42])  );
    wire logic pp_15_43;
    assign pp_15_43 = (select_e_15 & IN2[43] | select_2x_15 & IN2[42] | select_n2x_15 & (~ IN2[42]) | select_ne_15 & (~ IN2[43])  );
    wire logic pp_15_44;
    assign pp_15_44 = (select_e_15 & IN2[44] | select_2x_15 & IN2[43] | select_n2x_15 & (~ IN2[43]) | select_ne_15 & (~ IN2[44])  );
    wire logic pp_15_45;
    assign pp_15_45 = (select_e_15 & IN2[45] | select_2x_15 & IN2[44] | select_n2x_15 & (~ IN2[44]) | select_ne_15 & (~ IN2[45])  );
    wire logic pp_15_46;
    assign pp_15_46 = (select_e_15 & IN2[46] | select_2x_15 & IN2[45] | select_n2x_15 & (~ IN2[45]) | select_ne_15 & (~ IN2[46])  );
    wire logic pp_15_47;
    assign pp_15_47 = (select_e_15 & IN2[47] | select_2x_15 & IN2[46] | select_n2x_15 & (~ IN2[46]) | select_ne_15 & (~ IN2[47])  );
    wire logic pp_15_48;
    assign pp_15_48 = (select_e_15 & IN2[48] | select_2x_15 & IN2[47] | select_n2x_15 & (~ IN2[47]) | select_ne_15 & (~ IN2[48])  );
    wire logic pp_15_49;
    assign pp_15_49 = (select_e_15 & IN2[49] | select_2x_15 & IN2[48] | select_n2x_15 & (~ IN2[48]) | select_ne_15 & (~ IN2[49])  );
    wire logic pp_15_50;
    assign pp_15_50 = (select_e_15 & IN2[50] | select_2x_15 & IN2[49] | select_n2x_15 & (~ IN2[49]) | select_ne_15 & (~ IN2[50])  );
    wire logic pp_15_51;
    assign pp_15_51 = (select_e_15 & IN2[51] | select_2x_15 & IN2[50] | select_n2x_15 & (~ IN2[50]) | select_ne_15 & (~ IN2[51])  );
    wire logic pp_15_52;
    assign pp_15_52 = (select_e_15 & IN2[52] | select_2x_15 & IN2[51] | select_n2x_15 & (~ IN2[51]) | select_ne_15 & (~ IN2[52])  );
    wire logic pp_15_53;
    assign pp_15_53 = (select_e_15 & IN2[53] | select_2x_15 & IN2[52] | select_n2x_15 & (~ IN2[52]) | select_ne_15 & (~ IN2[53])  );
    wire logic pp_15_54;
    assign pp_15_54 = (select_e_15 & IN2[54] | select_2x_15 & IN2[53] | select_n2x_15 & (~ IN2[53]) | select_ne_15 & (~ IN2[54])  );
    wire logic pp_15_55;
    assign pp_15_55 = (select_e_15 & IN2[55] | select_2x_15 & IN2[54] | select_n2x_15 & (~ IN2[54]) | select_ne_15 & (~ IN2[55])  );
    wire logic pp_15_56;
    assign pp_15_56 = (select_e_15 & IN2[56] | select_2x_15 & IN2[55] | select_n2x_15 & (~ IN2[55]) | select_ne_15 & (~ IN2[56])  );
    wire logic pp_15_57;
    assign pp_15_57 = (select_e_15 & IN2[57] | select_2x_15 & IN2[56] | select_n2x_15 & (~ IN2[56]) | select_ne_15 & (~ IN2[57])  );
    wire logic pp_15_58;
    assign pp_15_58 = (select_e_15 & IN2[58] | select_2x_15 & IN2[57] | select_n2x_15 & (~ IN2[57]) | select_ne_15 & (~ IN2[58])  );
    wire logic pp_15_59;
    assign pp_15_59 = (select_e_15 & IN2[59] | select_2x_15 & IN2[58] | select_n2x_15 & (~ IN2[58]) | select_ne_15 & (~ IN2[59])  );
    wire logic pp_15_60;
    assign pp_15_60 = (select_e_15 & IN2[60] | select_2x_15 & IN2[59] | select_n2x_15 & (~ IN2[59]) | select_ne_15 & (~ IN2[60])  );
    wire logic pp_15_61;
    assign pp_15_61 = (select_e_15 & IN2[61] | select_2x_15 & IN2[60] | select_n2x_15 & (~ IN2[60]) | select_ne_15 & (~ IN2[61])  );
    wire logic pp_15_62;
    assign pp_15_62 = (select_e_15 & IN2[62] | select_2x_15 & IN2[61] | select_n2x_15 & (~ IN2[61]) | select_ne_15 & (~ IN2[62])  );
    wire logic pp_15_63;
    assign pp_15_63 = (select_e_15 & IN2[63] | select_2x_15 & IN2[62] | select_n2x_15 & (~ IN2[62]) | select_ne_15 & (~ IN2[63])  );
    wire logic pp_15_64;
    assign pp_15_64 = (select_e_15 & IN2[63] | select_2x_15 & IN2[63] | select_n2x_15 & (~ IN2[63]) | select_ne_15 & (~ IN2[63])  );
    wire logic pp_15_65;
    assign pp_15_65 = ~ (select_e_15 & IN2[63] | select_2x_15 & IN2[63] | select_n2x_15 & (~ IN2[63]) | select_ne_15 & (~ IN2[63])  );
    assign tcomp15 = select_ne_15 | select_n2x_15;
    
    // Signed Booth Radix-4 Partial Products Row 17
    wire logic select_e_16, select_ne_16, select_2x_16, tcomp16, select_n2x_16;
    assign select_e_16 = ((~ IN1[33]) & (IN1[32] ^ IN1[31]));
    assign select_ne_16 = IN1[33] &  (IN1[32] ^ IN1[31]);
    assign select_2x_16 = (~ IN1[33]) & IN1[32] & IN1[31];
    assign select_n2x_16 = IN1[33] & (~ IN1[32]) & (~ IN1[31]);
    wire logic pp_16_0;
    assign pp_16_0 = (select_e_16 & IN2[0] | select_2x_16 & 1'b0 | select_n2x_16 & 1'b1 | select_ne_16 & (~ IN2[0])  );
    wire logic pp_16_1;
    assign pp_16_1 = (select_e_16 & IN2[1] | select_2x_16 & IN2[0] | select_n2x_16 & (~ IN2[0]) | select_ne_16 & (~ IN2[1])  );
    wire logic pp_16_2;
    assign pp_16_2 = (select_e_16 & IN2[2] | select_2x_16 & IN2[1] | select_n2x_16 & (~ IN2[1]) | select_ne_16 & (~ IN2[2])  );
    wire logic pp_16_3;
    assign pp_16_3 = (select_e_16 & IN2[3] | select_2x_16 & IN2[2] | select_n2x_16 & (~ IN2[2]) | select_ne_16 & (~ IN2[3])  );
    wire logic pp_16_4;
    assign pp_16_4 = (select_e_16 & IN2[4] | select_2x_16 & IN2[3] | select_n2x_16 & (~ IN2[3]) | select_ne_16 & (~ IN2[4])  );
    wire logic pp_16_5;
    assign pp_16_5 = (select_e_16 & IN2[5] | select_2x_16 & IN2[4] | select_n2x_16 & (~ IN2[4]) | select_ne_16 & (~ IN2[5])  );
    wire logic pp_16_6;
    assign pp_16_6 = (select_e_16 & IN2[6] | select_2x_16 & IN2[5] | select_n2x_16 & (~ IN2[5]) | select_ne_16 & (~ IN2[6])  );
    wire logic pp_16_7;
    assign pp_16_7 = (select_e_16 & IN2[7] | select_2x_16 & IN2[6] | select_n2x_16 & (~ IN2[6]) | select_ne_16 & (~ IN2[7])  );
    wire logic pp_16_8;
    assign pp_16_8 = (select_e_16 & IN2[8] | select_2x_16 & IN2[7] | select_n2x_16 & (~ IN2[7]) | select_ne_16 & (~ IN2[8])  );
    wire logic pp_16_9;
    assign pp_16_9 = (select_e_16 & IN2[9] | select_2x_16 & IN2[8] | select_n2x_16 & (~ IN2[8]) | select_ne_16 & (~ IN2[9])  );
    wire logic pp_16_10;
    assign pp_16_10 = (select_e_16 & IN2[10] | select_2x_16 & IN2[9] | select_n2x_16 & (~ IN2[9]) | select_ne_16 & (~ IN2[10])  );
    wire logic pp_16_11;
    assign pp_16_11 = (select_e_16 & IN2[11] | select_2x_16 & IN2[10] | select_n2x_16 & (~ IN2[10]) | select_ne_16 & (~ IN2[11])  );
    wire logic pp_16_12;
    assign pp_16_12 = (select_e_16 & IN2[12] | select_2x_16 & IN2[11] | select_n2x_16 & (~ IN2[11]) | select_ne_16 & (~ IN2[12])  );
    wire logic pp_16_13;
    assign pp_16_13 = (select_e_16 & IN2[13] | select_2x_16 & IN2[12] | select_n2x_16 & (~ IN2[12]) | select_ne_16 & (~ IN2[13])  );
    wire logic pp_16_14;
    assign pp_16_14 = (select_e_16 & IN2[14] | select_2x_16 & IN2[13] | select_n2x_16 & (~ IN2[13]) | select_ne_16 & (~ IN2[14])  );
    wire logic pp_16_15;
    assign pp_16_15 = (select_e_16 & IN2[15] | select_2x_16 & IN2[14] | select_n2x_16 & (~ IN2[14]) | select_ne_16 & (~ IN2[15])  );
    wire logic pp_16_16;
    assign pp_16_16 = (select_e_16 & IN2[16] | select_2x_16 & IN2[15] | select_n2x_16 & (~ IN2[15]) | select_ne_16 & (~ IN2[16])  );
    wire logic pp_16_17;
    assign pp_16_17 = (select_e_16 & IN2[17] | select_2x_16 & IN2[16] | select_n2x_16 & (~ IN2[16]) | select_ne_16 & (~ IN2[17])  );
    wire logic pp_16_18;
    assign pp_16_18 = (select_e_16 & IN2[18] | select_2x_16 & IN2[17] | select_n2x_16 & (~ IN2[17]) | select_ne_16 & (~ IN2[18])  );
    wire logic pp_16_19;
    assign pp_16_19 = (select_e_16 & IN2[19] | select_2x_16 & IN2[18] | select_n2x_16 & (~ IN2[18]) | select_ne_16 & (~ IN2[19])  );
    wire logic pp_16_20;
    assign pp_16_20 = (select_e_16 & IN2[20] | select_2x_16 & IN2[19] | select_n2x_16 & (~ IN2[19]) | select_ne_16 & (~ IN2[20])  );
    wire logic pp_16_21;
    assign pp_16_21 = (select_e_16 & IN2[21] | select_2x_16 & IN2[20] | select_n2x_16 & (~ IN2[20]) | select_ne_16 & (~ IN2[21])  );
    wire logic pp_16_22;
    assign pp_16_22 = (select_e_16 & IN2[22] | select_2x_16 & IN2[21] | select_n2x_16 & (~ IN2[21]) | select_ne_16 & (~ IN2[22])  );
    wire logic pp_16_23;
    assign pp_16_23 = (select_e_16 & IN2[23] | select_2x_16 & IN2[22] | select_n2x_16 & (~ IN2[22]) | select_ne_16 & (~ IN2[23])  );
    wire logic pp_16_24;
    assign pp_16_24 = (select_e_16 & IN2[24] | select_2x_16 & IN2[23] | select_n2x_16 & (~ IN2[23]) | select_ne_16 & (~ IN2[24])  );
    wire logic pp_16_25;
    assign pp_16_25 = (select_e_16 & IN2[25] | select_2x_16 & IN2[24] | select_n2x_16 & (~ IN2[24]) | select_ne_16 & (~ IN2[25])  );
    wire logic pp_16_26;
    assign pp_16_26 = (select_e_16 & IN2[26] | select_2x_16 & IN2[25] | select_n2x_16 & (~ IN2[25]) | select_ne_16 & (~ IN2[26])  );
    wire logic pp_16_27;
    assign pp_16_27 = (select_e_16 & IN2[27] | select_2x_16 & IN2[26] | select_n2x_16 & (~ IN2[26]) | select_ne_16 & (~ IN2[27])  );
    wire logic pp_16_28;
    assign pp_16_28 = (select_e_16 & IN2[28] | select_2x_16 & IN2[27] | select_n2x_16 & (~ IN2[27]) | select_ne_16 & (~ IN2[28])  );
    wire logic pp_16_29;
    assign pp_16_29 = (select_e_16 & IN2[29] | select_2x_16 & IN2[28] | select_n2x_16 & (~ IN2[28]) | select_ne_16 & (~ IN2[29])  );
    wire logic pp_16_30;
    assign pp_16_30 = (select_e_16 & IN2[30] | select_2x_16 & IN2[29] | select_n2x_16 & (~ IN2[29]) | select_ne_16 & (~ IN2[30])  );
    wire logic pp_16_31;
    assign pp_16_31 = (select_e_16 & IN2[31] | select_2x_16 & IN2[30] | select_n2x_16 & (~ IN2[30]) | select_ne_16 & (~ IN2[31])  );
    wire logic pp_16_32;
    assign pp_16_32 = (select_e_16 & IN2[32] | select_2x_16 & IN2[31] | select_n2x_16 & (~ IN2[31]) | select_ne_16 & (~ IN2[32])  );
    wire logic pp_16_33;
    assign pp_16_33 = (select_e_16 & IN2[33] | select_2x_16 & IN2[32] | select_n2x_16 & (~ IN2[32]) | select_ne_16 & (~ IN2[33])  );
    wire logic pp_16_34;
    assign pp_16_34 = (select_e_16 & IN2[34] | select_2x_16 & IN2[33] | select_n2x_16 & (~ IN2[33]) | select_ne_16 & (~ IN2[34])  );
    wire logic pp_16_35;
    assign pp_16_35 = (select_e_16 & IN2[35] | select_2x_16 & IN2[34] | select_n2x_16 & (~ IN2[34]) | select_ne_16 & (~ IN2[35])  );
    wire logic pp_16_36;
    assign pp_16_36 = (select_e_16 & IN2[36] | select_2x_16 & IN2[35] | select_n2x_16 & (~ IN2[35]) | select_ne_16 & (~ IN2[36])  );
    wire logic pp_16_37;
    assign pp_16_37 = (select_e_16 & IN2[37] | select_2x_16 & IN2[36] | select_n2x_16 & (~ IN2[36]) | select_ne_16 & (~ IN2[37])  );
    wire logic pp_16_38;
    assign pp_16_38 = (select_e_16 & IN2[38] | select_2x_16 & IN2[37] | select_n2x_16 & (~ IN2[37]) | select_ne_16 & (~ IN2[38])  );
    wire logic pp_16_39;
    assign pp_16_39 = (select_e_16 & IN2[39] | select_2x_16 & IN2[38] | select_n2x_16 & (~ IN2[38]) | select_ne_16 & (~ IN2[39])  );
    wire logic pp_16_40;
    assign pp_16_40 = (select_e_16 & IN2[40] | select_2x_16 & IN2[39] | select_n2x_16 & (~ IN2[39]) | select_ne_16 & (~ IN2[40])  );
    wire logic pp_16_41;
    assign pp_16_41 = (select_e_16 & IN2[41] | select_2x_16 & IN2[40] | select_n2x_16 & (~ IN2[40]) | select_ne_16 & (~ IN2[41])  );
    wire logic pp_16_42;
    assign pp_16_42 = (select_e_16 & IN2[42] | select_2x_16 & IN2[41] | select_n2x_16 & (~ IN2[41]) | select_ne_16 & (~ IN2[42])  );
    wire logic pp_16_43;
    assign pp_16_43 = (select_e_16 & IN2[43] | select_2x_16 & IN2[42] | select_n2x_16 & (~ IN2[42]) | select_ne_16 & (~ IN2[43])  );
    wire logic pp_16_44;
    assign pp_16_44 = (select_e_16 & IN2[44] | select_2x_16 & IN2[43] | select_n2x_16 & (~ IN2[43]) | select_ne_16 & (~ IN2[44])  );
    wire logic pp_16_45;
    assign pp_16_45 = (select_e_16 & IN2[45] | select_2x_16 & IN2[44] | select_n2x_16 & (~ IN2[44]) | select_ne_16 & (~ IN2[45])  );
    wire logic pp_16_46;
    assign pp_16_46 = (select_e_16 & IN2[46] | select_2x_16 & IN2[45] | select_n2x_16 & (~ IN2[45]) | select_ne_16 & (~ IN2[46])  );
    wire logic pp_16_47;
    assign pp_16_47 = (select_e_16 & IN2[47] | select_2x_16 & IN2[46] | select_n2x_16 & (~ IN2[46]) | select_ne_16 & (~ IN2[47])  );
    wire logic pp_16_48;
    assign pp_16_48 = (select_e_16 & IN2[48] | select_2x_16 & IN2[47] | select_n2x_16 & (~ IN2[47]) | select_ne_16 & (~ IN2[48])  );
    wire logic pp_16_49;
    assign pp_16_49 = (select_e_16 & IN2[49] | select_2x_16 & IN2[48] | select_n2x_16 & (~ IN2[48]) | select_ne_16 & (~ IN2[49])  );
    wire logic pp_16_50;
    assign pp_16_50 = (select_e_16 & IN2[50] | select_2x_16 & IN2[49] | select_n2x_16 & (~ IN2[49]) | select_ne_16 & (~ IN2[50])  );
    wire logic pp_16_51;
    assign pp_16_51 = (select_e_16 & IN2[51] | select_2x_16 & IN2[50] | select_n2x_16 & (~ IN2[50]) | select_ne_16 & (~ IN2[51])  );
    wire logic pp_16_52;
    assign pp_16_52 = (select_e_16 & IN2[52] | select_2x_16 & IN2[51] | select_n2x_16 & (~ IN2[51]) | select_ne_16 & (~ IN2[52])  );
    wire logic pp_16_53;
    assign pp_16_53 = (select_e_16 & IN2[53] | select_2x_16 & IN2[52] | select_n2x_16 & (~ IN2[52]) | select_ne_16 & (~ IN2[53])  );
    wire logic pp_16_54;
    assign pp_16_54 = (select_e_16 & IN2[54] | select_2x_16 & IN2[53] | select_n2x_16 & (~ IN2[53]) | select_ne_16 & (~ IN2[54])  );
    wire logic pp_16_55;
    assign pp_16_55 = (select_e_16 & IN2[55] | select_2x_16 & IN2[54] | select_n2x_16 & (~ IN2[54]) | select_ne_16 & (~ IN2[55])  );
    wire logic pp_16_56;
    assign pp_16_56 = (select_e_16 & IN2[56] | select_2x_16 & IN2[55] | select_n2x_16 & (~ IN2[55]) | select_ne_16 & (~ IN2[56])  );
    wire logic pp_16_57;
    assign pp_16_57 = (select_e_16 & IN2[57] | select_2x_16 & IN2[56] | select_n2x_16 & (~ IN2[56]) | select_ne_16 & (~ IN2[57])  );
    wire logic pp_16_58;
    assign pp_16_58 = (select_e_16 & IN2[58] | select_2x_16 & IN2[57] | select_n2x_16 & (~ IN2[57]) | select_ne_16 & (~ IN2[58])  );
    wire logic pp_16_59;
    assign pp_16_59 = (select_e_16 & IN2[59] | select_2x_16 & IN2[58] | select_n2x_16 & (~ IN2[58]) | select_ne_16 & (~ IN2[59])  );
    wire logic pp_16_60;
    assign pp_16_60 = (select_e_16 & IN2[60] | select_2x_16 & IN2[59] | select_n2x_16 & (~ IN2[59]) | select_ne_16 & (~ IN2[60])  );
    wire logic pp_16_61;
    assign pp_16_61 = (select_e_16 & IN2[61] | select_2x_16 & IN2[60] | select_n2x_16 & (~ IN2[60]) | select_ne_16 & (~ IN2[61])  );
    wire logic pp_16_62;
    assign pp_16_62 = (select_e_16 & IN2[62] | select_2x_16 & IN2[61] | select_n2x_16 & (~ IN2[61]) | select_ne_16 & (~ IN2[62])  );
    wire logic pp_16_63;
    assign pp_16_63 = (select_e_16 & IN2[63] | select_2x_16 & IN2[62] | select_n2x_16 & (~ IN2[62]) | select_ne_16 & (~ IN2[63])  );
    wire logic pp_16_64;
    assign pp_16_64 = (select_e_16 & IN2[63] | select_2x_16 & IN2[63] | select_n2x_16 & (~ IN2[63]) | select_ne_16 & (~ IN2[63])  );
    wire logic pp_16_65;
    assign pp_16_65 = ~ (select_e_16 & IN2[63] | select_2x_16 & IN2[63] | select_n2x_16 & (~ IN2[63]) | select_ne_16 & (~ IN2[63])  );
    assign tcomp16 = select_ne_16 | select_n2x_16;
    
    // Signed Booth Radix-4 Partial Products Row 18
    wire logic select_e_17, select_ne_17, select_2x_17, tcomp17, select_n2x_17;
    assign select_e_17 = ((~ IN1[35]) & (IN1[34] ^ IN1[33]));
    assign select_ne_17 = IN1[35] &  (IN1[34] ^ IN1[33]);
    assign select_2x_17 = (~ IN1[35]) & IN1[34] & IN1[33];
    assign select_n2x_17 = IN1[35] & (~ IN1[34]) & (~ IN1[33]);
    wire logic pp_17_0;
    assign pp_17_0 = (select_e_17 & IN2[0] | select_2x_17 & 1'b0 | select_n2x_17 & 1'b1 | select_ne_17 & (~ IN2[0])  );
    wire logic pp_17_1;
    assign pp_17_1 = (select_e_17 & IN2[1] | select_2x_17 & IN2[0] | select_n2x_17 & (~ IN2[0]) | select_ne_17 & (~ IN2[1])  );
    wire logic pp_17_2;
    assign pp_17_2 = (select_e_17 & IN2[2] | select_2x_17 & IN2[1] | select_n2x_17 & (~ IN2[1]) | select_ne_17 & (~ IN2[2])  );
    wire logic pp_17_3;
    assign pp_17_3 = (select_e_17 & IN2[3] | select_2x_17 & IN2[2] | select_n2x_17 & (~ IN2[2]) | select_ne_17 & (~ IN2[3])  );
    wire logic pp_17_4;
    assign pp_17_4 = (select_e_17 & IN2[4] | select_2x_17 & IN2[3] | select_n2x_17 & (~ IN2[3]) | select_ne_17 & (~ IN2[4])  );
    wire logic pp_17_5;
    assign pp_17_5 = (select_e_17 & IN2[5] | select_2x_17 & IN2[4] | select_n2x_17 & (~ IN2[4]) | select_ne_17 & (~ IN2[5])  );
    wire logic pp_17_6;
    assign pp_17_6 = (select_e_17 & IN2[6] | select_2x_17 & IN2[5] | select_n2x_17 & (~ IN2[5]) | select_ne_17 & (~ IN2[6])  );
    wire logic pp_17_7;
    assign pp_17_7 = (select_e_17 & IN2[7] | select_2x_17 & IN2[6] | select_n2x_17 & (~ IN2[6]) | select_ne_17 & (~ IN2[7])  );
    wire logic pp_17_8;
    assign pp_17_8 = (select_e_17 & IN2[8] | select_2x_17 & IN2[7] | select_n2x_17 & (~ IN2[7]) | select_ne_17 & (~ IN2[8])  );
    wire logic pp_17_9;
    assign pp_17_9 = (select_e_17 & IN2[9] | select_2x_17 & IN2[8] | select_n2x_17 & (~ IN2[8]) | select_ne_17 & (~ IN2[9])  );
    wire logic pp_17_10;
    assign pp_17_10 = (select_e_17 & IN2[10] | select_2x_17 & IN2[9] | select_n2x_17 & (~ IN2[9]) | select_ne_17 & (~ IN2[10])  );
    wire logic pp_17_11;
    assign pp_17_11 = (select_e_17 & IN2[11] | select_2x_17 & IN2[10] | select_n2x_17 & (~ IN2[10]) | select_ne_17 & (~ IN2[11])  );
    wire logic pp_17_12;
    assign pp_17_12 = (select_e_17 & IN2[12] | select_2x_17 & IN2[11] | select_n2x_17 & (~ IN2[11]) | select_ne_17 & (~ IN2[12])  );
    wire logic pp_17_13;
    assign pp_17_13 = (select_e_17 & IN2[13] | select_2x_17 & IN2[12] | select_n2x_17 & (~ IN2[12]) | select_ne_17 & (~ IN2[13])  );
    wire logic pp_17_14;
    assign pp_17_14 = (select_e_17 & IN2[14] | select_2x_17 & IN2[13] | select_n2x_17 & (~ IN2[13]) | select_ne_17 & (~ IN2[14])  );
    wire logic pp_17_15;
    assign pp_17_15 = (select_e_17 & IN2[15] | select_2x_17 & IN2[14] | select_n2x_17 & (~ IN2[14]) | select_ne_17 & (~ IN2[15])  );
    wire logic pp_17_16;
    assign pp_17_16 = (select_e_17 & IN2[16] | select_2x_17 & IN2[15] | select_n2x_17 & (~ IN2[15]) | select_ne_17 & (~ IN2[16])  );
    wire logic pp_17_17;
    assign pp_17_17 = (select_e_17 & IN2[17] | select_2x_17 & IN2[16] | select_n2x_17 & (~ IN2[16]) | select_ne_17 & (~ IN2[17])  );
    wire logic pp_17_18;
    assign pp_17_18 = (select_e_17 & IN2[18] | select_2x_17 & IN2[17] | select_n2x_17 & (~ IN2[17]) | select_ne_17 & (~ IN2[18])  );
    wire logic pp_17_19;
    assign pp_17_19 = (select_e_17 & IN2[19] | select_2x_17 & IN2[18] | select_n2x_17 & (~ IN2[18]) | select_ne_17 & (~ IN2[19])  );
    wire logic pp_17_20;
    assign pp_17_20 = (select_e_17 & IN2[20] | select_2x_17 & IN2[19] | select_n2x_17 & (~ IN2[19]) | select_ne_17 & (~ IN2[20])  );
    wire logic pp_17_21;
    assign pp_17_21 = (select_e_17 & IN2[21] | select_2x_17 & IN2[20] | select_n2x_17 & (~ IN2[20]) | select_ne_17 & (~ IN2[21])  );
    wire logic pp_17_22;
    assign pp_17_22 = (select_e_17 & IN2[22] | select_2x_17 & IN2[21] | select_n2x_17 & (~ IN2[21]) | select_ne_17 & (~ IN2[22])  );
    wire logic pp_17_23;
    assign pp_17_23 = (select_e_17 & IN2[23] | select_2x_17 & IN2[22] | select_n2x_17 & (~ IN2[22]) | select_ne_17 & (~ IN2[23])  );
    wire logic pp_17_24;
    assign pp_17_24 = (select_e_17 & IN2[24] | select_2x_17 & IN2[23] | select_n2x_17 & (~ IN2[23]) | select_ne_17 & (~ IN2[24])  );
    wire logic pp_17_25;
    assign pp_17_25 = (select_e_17 & IN2[25] | select_2x_17 & IN2[24] | select_n2x_17 & (~ IN2[24]) | select_ne_17 & (~ IN2[25])  );
    wire logic pp_17_26;
    assign pp_17_26 = (select_e_17 & IN2[26] | select_2x_17 & IN2[25] | select_n2x_17 & (~ IN2[25]) | select_ne_17 & (~ IN2[26])  );
    wire logic pp_17_27;
    assign pp_17_27 = (select_e_17 & IN2[27] | select_2x_17 & IN2[26] | select_n2x_17 & (~ IN2[26]) | select_ne_17 & (~ IN2[27])  );
    wire logic pp_17_28;
    assign pp_17_28 = (select_e_17 & IN2[28] | select_2x_17 & IN2[27] | select_n2x_17 & (~ IN2[27]) | select_ne_17 & (~ IN2[28])  );
    wire logic pp_17_29;
    assign pp_17_29 = (select_e_17 & IN2[29] | select_2x_17 & IN2[28] | select_n2x_17 & (~ IN2[28]) | select_ne_17 & (~ IN2[29])  );
    wire logic pp_17_30;
    assign pp_17_30 = (select_e_17 & IN2[30] | select_2x_17 & IN2[29] | select_n2x_17 & (~ IN2[29]) | select_ne_17 & (~ IN2[30])  );
    wire logic pp_17_31;
    assign pp_17_31 = (select_e_17 & IN2[31] | select_2x_17 & IN2[30] | select_n2x_17 & (~ IN2[30]) | select_ne_17 & (~ IN2[31])  );
    wire logic pp_17_32;
    assign pp_17_32 = (select_e_17 & IN2[32] | select_2x_17 & IN2[31] | select_n2x_17 & (~ IN2[31]) | select_ne_17 & (~ IN2[32])  );
    wire logic pp_17_33;
    assign pp_17_33 = (select_e_17 & IN2[33] | select_2x_17 & IN2[32] | select_n2x_17 & (~ IN2[32]) | select_ne_17 & (~ IN2[33])  );
    wire logic pp_17_34;
    assign pp_17_34 = (select_e_17 & IN2[34] | select_2x_17 & IN2[33] | select_n2x_17 & (~ IN2[33]) | select_ne_17 & (~ IN2[34])  );
    wire logic pp_17_35;
    assign pp_17_35 = (select_e_17 & IN2[35] | select_2x_17 & IN2[34] | select_n2x_17 & (~ IN2[34]) | select_ne_17 & (~ IN2[35])  );
    wire logic pp_17_36;
    assign pp_17_36 = (select_e_17 & IN2[36] | select_2x_17 & IN2[35] | select_n2x_17 & (~ IN2[35]) | select_ne_17 & (~ IN2[36])  );
    wire logic pp_17_37;
    assign pp_17_37 = (select_e_17 & IN2[37] | select_2x_17 & IN2[36] | select_n2x_17 & (~ IN2[36]) | select_ne_17 & (~ IN2[37])  );
    wire logic pp_17_38;
    assign pp_17_38 = (select_e_17 & IN2[38] | select_2x_17 & IN2[37] | select_n2x_17 & (~ IN2[37]) | select_ne_17 & (~ IN2[38])  );
    wire logic pp_17_39;
    assign pp_17_39 = (select_e_17 & IN2[39] | select_2x_17 & IN2[38] | select_n2x_17 & (~ IN2[38]) | select_ne_17 & (~ IN2[39])  );
    wire logic pp_17_40;
    assign pp_17_40 = (select_e_17 & IN2[40] | select_2x_17 & IN2[39] | select_n2x_17 & (~ IN2[39]) | select_ne_17 & (~ IN2[40])  );
    wire logic pp_17_41;
    assign pp_17_41 = (select_e_17 & IN2[41] | select_2x_17 & IN2[40] | select_n2x_17 & (~ IN2[40]) | select_ne_17 & (~ IN2[41])  );
    wire logic pp_17_42;
    assign pp_17_42 = (select_e_17 & IN2[42] | select_2x_17 & IN2[41] | select_n2x_17 & (~ IN2[41]) | select_ne_17 & (~ IN2[42])  );
    wire logic pp_17_43;
    assign pp_17_43 = (select_e_17 & IN2[43] | select_2x_17 & IN2[42] | select_n2x_17 & (~ IN2[42]) | select_ne_17 & (~ IN2[43])  );
    wire logic pp_17_44;
    assign pp_17_44 = (select_e_17 & IN2[44] | select_2x_17 & IN2[43] | select_n2x_17 & (~ IN2[43]) | select_ne_17 & (~ IN2[44])  );
    wire logic pp_17_45;
    assign pp_17_45 = (select_e_17 & IN2[45] | select_2x_17 & IN2[44] | select_n2x_17 & (~ IN2[44]) | select_ne_17 & (~ IN2[45])  );
    wire logic pp_17_46;
    assign pp_17_46 = (select_e_17 & IN2[46] | select_2x_17 & IN2[45] | select_n2x_17 & (~ IN2[45]) | select_ne_17 & (~ IN2[46])  );
    wire logic pp_17_47;
    assign pp_17_47 = (select_e_17 & IN2[47] | select_2x_17 & IN2[46] | select_n2x_17 & (~ IN2[46]) | select_ne_17 & (~ IN2[47])  );
    wire logic pp_17_48;
    assign pp_17_48 = (select_e_17 & IN2[48] | select_2x_17 & IN2[47] | select_n2x_17 & (~ IN2[47]) | select_ne_17 & (~ IN2[48])  );
    wire logic pp_17_49;
    assign pp_17_49 = (select_e_17 & IN2[49] | select_2x_17 & IN2[48] | select_n2x_17 & (~ IN2[48]) | select_ne_17 & (~ IN2[49])  );
    wire logic pp_17_50;
    assign pp_17_50 = (select_e_17 & IN2[50] | select_2x_17 & IN2[49] | select_n2x_17 & (~ IN2[49]) | select_ne_17 & (~ IN2[50])  );
    wire logic pp_17_51;
    assign pp_17_51 = (select_e_17 & IN2[51] | select_2x_17 & IN2[50] | select_n2x_17 & (~ IN2[50]) | select_ne_17 & (~ IN2[51])  );
    wire logic pp_17_52;
    assign pp_17_52 = (select_e_17 & IN2[52] | select_2x_17 & IN2[51] | select_n2x_17 & (~ IN2[51]) | select_ne_17 & (~ IN2[52])  );
    wire logic pp_17_53;
    assign pp_17_53 = (select_e_17 & IN2[53] | select_2x_17 & IN2[52] | select_n2x_17 & (~ IN2[52]) | select_ne_17 & (~ IN2[53])  );
    wire logic pp_17_54;
    assign pp_17_54 = (select_e_17 & IN2[54] | select_2x_17 & IN2[53] | select_n2x_17 & (~ IN2[53]) | select_ne_17 & (~ IN2[54])  );
    wire logic pp_17_55;
    assign pp_17_55 = (select_e_17 & IN2[55] | select_2x_17 & IN2[54] | select_n2x_17 & (~ IN2[54]) | select_ne_17 & (~ IN2[55])  );
    wire logic pp_17_56;
    assign pp_17_56 = (select_e_17 & IN2[56] | select_2x_17 & IN2[55] | select_n2x_17 & (~ IN2[55]) | select_ne_17 & (~ IN2[56])  );
    wire logic pp_17_57;
    assign pp_17_57 = (select_e_17 & IN2[57] | select_2x_17 & IN2[56] | select_n2x_17 & (~ IN2[56]) | select_ne_17 & (~ IN2[57])  );
    wire logic pp_17_58;
    assign pp_17_58 = (select_e_17 & IN2[58] | select_2x_17 & IN2[57] | select_n2x_17 & (~ IN2[57]) | select_ne_17 & (~ IN2[58])  );
    wire logic pp_17_59;
    assign pp_17_59 = (select_e_17 & IN2[59] | select_2x_17 & IN2[58] | select_n2x_17 & (~ IN2[58]) | select_ne_17 & (~ IN2[59])  );
    wire logic pp_17_60;
    assign pp_17_60 = (select_e_17 & IN2[60] | select_2x_17 & IN2[59] | select_n2x_17 & (~ IN2[59]) | select_ne_17 & (~ IN2[60])  );
    wire logic pp_17_61;
    assign pp_17_61 = (select_e_17 & IN2[61] | select_2x_17 & IN2[60] | select_n2x_17 & (~ IN2[60]) | select_ne_17 & (~ IN2[61])  );
    wire logic pp_17_62;
    assign pp_17_62 = (select_e_17 & IN2[62] | select_2x_17 & IN2[61] | select_n2x_17 & (~ IN2[61]) | select_ne_17 & (~ IN2[62])  );
    wire logic pp_17_63;
    assign pp_17_63 = (select_e_17 & IN2[63] | select_2x_17 & IN2[62] | select_n2x_17 & (~ IN2[62]) | select_ne_17 & (~ IN2[63])  );
    wire logic pp_17_64;
    assign pp_17_64 = (select_e_17 & IN2[63] | select_2x_17 & IN2[63] | select_n2x_17 & (~ IN2[63]) | select_ne_17 & (~ IN2[63])  );
    wire logic pp_17_65;
    assign pp_17_65 = ~ (select_e_17 & IN2[63] | select_2x_17 & IN2[63] | select_n2x_17 & (~ IN2[63]) | select_ne_17 & (~ IN2[63])  );
    assign tcomp17 = select_ne_17 | select_n2x_17;
    
    // Signed Booth Radix-4 Partial Products Row 19
    wire logic select_e_18, select_ne_18, select_2x_18, tcomp18, select_n2x_18;
    assign select_e_18 = ((~ IN1[37]) & (IN1[36] ^ IN1[35]));
    assign select_ne_18 = IN1[37] &  (IN1[36] ^ IN1[35]);
    assign select_2x_18 = (~ IN1[37]) & IN1[36] & IN1[35];
    assign select_n2x_18 = IN1[37] & (~ IN1[36]) & (~ IN1[35]);
    wire logic pp_18_0;
    assign pp_18_0 = (select_e_18 & IN2[0] | select_2x_18 & 1'b0 | select_n2x_18 & 1'b1 | select_ne_18 & (~ IN2[0])  );
    wire logic pp_18_1;
    assign pp_18_1 = (select_e_18 & IN2[1] | select_2x_18 & IN2[0] | select_n2x_18 & (~ IN2[0]) | select_ne_18 & (~ IN2[1])  );
    wire logic pp_18_2;
    assign pp_18_2 = (select_e_18 & IN2[2] | select_2x_18 & IN2[1] | select_n2x_18 & (~ IN2[1]) | select_ne_18 & (~ IN2[2])  );
    wire logic pp_18_3;
    assign pp_18_3 = (select_e_18 & IN2[3] | select_2x_18 & IN2[2] | select_n2x_18 & (~ IN2[2]) | select_ne_18 & (~ IN2[3])  );
    wire logic pp_18_4;
    assign pp_18_4 = (select_e_18 & IN2[4] | select_2x_18 & IN2[3] | select_n2x_18 & (~ IN2[3]) | select_ne_18 & (~ IN2[4])  );
    wire logic pp_18_5;
    assign pp_18_5 = (select_e_18 & IN2[5] | select_2x_18 & IN2[4] | select_n2x_18 & (~ IN2[4]) | select_ne_18 & (~ IN2[5])  );
    wire logic pp_18_6;
    assign pp_18_6 = (select_e_18 & IN2[6] | select_2x_18 & IN2[5] | select_n2x_18 & (~ IN2[5]) | select_ne_18 & (~ IN2[6])  );
    wire logic pp_18_7;
    assign pp_18_7 = (select_e_18 & IN2[7] | select_2x_18 & IN2[6] | select_n2x_18 & (~ IN2[6]) | select_ne_18 & (~ IN2[7])  );
    wire logic pp_18_8;
    assign pp_18_8 = (select_e_18 & IN2[8] | select_2x_18 & IN2[7] | select_n2x_18 & (~ IN2[7]) | select_ne_18 & (~ IN2[8])  );
    wire logic pp_18_9;
    assign pp_18_9 = (select_e_18 & IN2[9] | select_2x_18 & IN2[8] | select_n2x_18 & (~ IN2[8]) | select_ne_18 & (~ IN2[9])  );
    wire logic pp_18_10;
    assign pp_18_10 = (select_e_18 & IN2[10] | select_2x_18 & IN2[9] | select_n2x_18 & (~ IN2[9]) | select_ne_18 & (~ IN2[10])  );
    wire logic pp_18_11;
    assign pp_18_11 = (select_e_18 & IN2[11] | select_2x_18 & IN2[10] | select_n2x_18 & (~ IN2[10]) | select_ne_18 & (~ IN2[11])  );
    wire logic pp_18_12;
    assign pp_18_12 = (select_e_18 & IN2[12] | select_2x_18 & IN2[11] | select_n2x_18 & (~ IN2[11]) | select_ne_18 & (~ IN2[12])  );
    wire logic pp_18_13;
    assign pp_18_13 = (select_e_18 & IN2[13] | select_2x_18 & IN2[12] | select_n2x_18 & (~ IN2[12]) | select_ne_18 & (~ IN2[13])  );
    wire logic pp_18_14;
    assign pp_18_14 = (select_e_18 & IN2[14] | select_2x_18 & IN2[13] | select_n2x_18 & (~ IN2[13]) | select_ne_18 & (~ IN2[14])  );
    wire logic pp_18_15;
    assign pp_18_15 = (select_e_18 & IN2[15] | select_2x_18 & IN2[14] | select_n2x_18 & (~ IN2[14]) | select_ne_18 & (~ IN2[15])  );
    wire logic pp_18_16;
    assign pp_18_16 = (select_e_18 & IN2[16] | select_2x_18 & IN2[15] | select_n2x_18 & (~ IN2[15]) | select_ne_18 & (~ IN2[16])  );
    wire logic pp_18_17;
    assign pp_18_17 = (select_e_18 & IN2[17] | select_2x_18 & IN2[16] | select_n2x_18 & (~ IN2[16]) | select_ne_18 & (~ IN2[17])  );
    wire logic pp_18_18;
    assign pp_18_18 = (select_e_18 & IN2[18] | select_2x_18 & IN2[17] | select_n2x_18 & (~ IN2[17]) | select_ne_18 & (~ IN2[18])  );
    wire logic pp_18_19;
    assign pp_18_19 = (select_e_18 & IN2[19] | select_2x_18 & IN2[18] | select_n2x_18 & (~ IN2[18]) | select_ne_18 & (~ IN2[19])  );
    wire logic pp_18_20;
    assign pp_18_20 = (select_e_18 & IN2[20] | select_2x_18 & IN2[19] | select_n2x_18 & (~ IN2[19]) | select_ne_18 & (~ IN2[20])  );
    wire logic pp_18_21;
    assign pp_18_21 = (select_e_18 & IN2[21] | select_2x_18 & IN2[20] | select_n2x_18 & (~ IN2[20]) | select_ne_18 & (~ IN2[21])  );
    wire logic pp_18_22;
    assign pp_18_22 = (select_e_18 & IN2[22] | select_2x_18 & IN2[21] | select_n2x_18 & (~ IN2[21]) | select_ne_18 & (~ IN2[22])  );
    wire logic pp_18_23;
    assign pp_18_23 = (select_e_18 & IN2[23] | select_2x_18 & IN2[22] | select_n2x_18 & (~ IN2[22]) | select_ne_18 & (~ IN2[23])  );
    wire logic pp_18_24;
    assign pp_18_24 = (select_e_18 & IN2[24] | select_2x_18 & IN2[23] | select_n2x_18 & (~ IN2[23]) | select_ne_18 & (~ IN2[24])  );
    wire logic pp_18_25;
    assign pp_18_25 = (select_e_18 & IN2[25] | select_2x_18 & IN2[24] | select_n2x_18 & (~ IN2[24]) | select_ne_18 & (~ IN2[25])  );
    wire logic pp_18_26;
    assign pp_18_26 = (select_e_18 & IN2[26] | select_2x_18 & IN2[25] | select_n2x_18 & (~ IN2[25]) | select_ne_18 & (~ IN2[26])  );
    wire logic pp_18_27;
    assign pp_18_27 = (select_e_18 & IN2[27] | select_2x_18 & IN2[26] | select_n2x_18 & (~ IN2[26]) | select_ne_18 & (~ IN2[27])  );
    wire logic pp_18_28;
    assign pp_18_28 = (select_e_18 & IN2[28] | select_2x_18 & IN2[27] | select_n2x_18 & (~ IN2[27]) | select_ne_18 & (~ IN2[28])  );
    wire logic pp_18_29;
    assign pp_18_29 = (select_e_18 & IN2[29] | select_2x_18 & IN2[28] | select_n2x_18 & (~ IN2[28]) | select_ne_18 & (~ IN2[29])  );
    wire logic pp_18_30;
    assign pp_18_30 = (select_e_18 & IN2[30] | select_2x_18 & IN2[29] | select_n2x_18 & (~ IN2[29]) | select_ne_18 & (~ IN2[30])  );
    wire logic pp_18_31;
    assign pp_18_31 = (select_e_18 & IN2[31] | select_2x_18 & IN2[30] | select_n2x_18 & (~ IN2[30]) | select_ne_18 & (~ IN2[31])  );
    wire logic pp_18_32;
    assign pp_18_32 = (select_e_18 & IN2[32] | select_2x_18 & IN2[31] | select_n2x_18 & (~ IN2[31]) | select_ne_18 & (~ IN2[32])  );
    wire logic pp_18_33;
    assign pp_18_33 = (select_e_18 & IN2[33] | select_2x_18 & IN2[32] | select_n2x_18 & (~ IN2[32]) | select_ne_18 & (~ IN2[33])  );
    wire logic pp_18_34;
    assign pp_18_34 = (select_e_18 & IN2[34] | select_2x_18 & IN2[33] | select_n2x_18 & (~ IN2[33]) | select_ne_18 & (~ IN2[34])  );
    wire logic pp_18_35;
    assign pp_18_35 = (select_e_18 & IN2[35] | select_2x_18 & IN2[34] | select_n2x_18 & (~ IN2[34]) | select_ne_18 & (~ IN2[35])  );
    wire logic pp_18_36;
    assign pp_18_36 = (select_e_18 & IN2[36] | select_2x_18 & IN2[35] | select_n2x_18 & (~ IN2[35]) | select_ne_18 & (~ IN2[36])  );
    wire logic pp_18_37;
    assign pp_18_37 = (select_e_18 & IN2[37] | select_2x_18 & IN2[36] | select_n2x_18 & (~ IN2[36]) | select_ne_18 & (~ IN2[37])  );
    wire logic pp_18_38;
    assign pp_18_38 = (select_e_18 & IN2[38] | select_2x_18 & IN2[37] | select_n2x_18 & (~ IN2[37]) | select_ne_18 & (~ IN2[38])  );
    wire logic pp_18_39;
    assign pp_18_39 = (select_e_18 & IN2[39] | select_2x_18 & IN2[38] | select_n2x_18 & (~ IN2[38]) | select_ne_18 & (~ IN2[39])  );
    wire logic pp_18_40;
    assign pp_18_40 = (select_e_18 & IN2[40] | select_2x_18 & IN2[39] | select_n2x_18 & (~ IN2[39]) | select_ne_18 & (~ IN2[40])  );
    wire logic pp_18_41;
    assign pp_18_41 = (select_e_18 & IN2[41] | select_2x_18 & IN2[40] | select_n2x_18 & (~ IN2[40]) | select_ne_18 & (~ IN2[41])  );
    wire logic pp_18_42;
    assign pp_18_42 = (select_e_18 & IN2[42] | select_2x_18 & IN2[41] | select_n2x_18 & (~ IN2[41]) | select_ne_18 & (~ IN2[42])  );
    wire logic pp_18_43;
    assign pp_18_43 = (select_e_18 & IN2[43] | select_2x_18 & IN2[42] | select_n2x_18 & (~ IN2[42]) | select_ne_18 & (~ IN2[43])  );
    wire logic pp_18_44;
    assign pp_18_44 = (select_e_18 & IN2[44] | select_2x_18 & IN2[43] | select_n2x_18 & (~ IN2[43]) | select_ne_18 & (~ IN2[44])  );
    wire logic pp_18_45;
    assign pp_18_45 = (select_e_18 & IN2[45] | select_2x_18 & IN2[44] | select_n2x_18 & (~ IN2[44]) | select_ne_18 & (~ IN2[45])  );
    wire logic pp_18_46;
    assign pp_18_46 = (select_e_18 & IN2[46] | select_2x_18 & IN2[45] | select_n2x_18 & (~ IN2[45]) | select_ne_18 & (~ IN2[46])  );
    wire logic pp_18_47;
    assign pp_18_47 = (select_e_18 & IN2[47] | select_2x_18 & IN2[46] | select_n2x_18 & (~ IN2[46]) | select_ne_18 & (~ IN2[47])  );
    wire logic pp_18_48;
    assign pp_18_48 = (select_e_18 & IN2[48] | select_2x_18 & IN2[47] | select_n2x_18 & (~ IN2[47]) | select_ne_18 & (~ IN2[48])  );
    wire logic pp_18_49;
    assign pp_18_49 = (select_e_18 & IN2[49] | select_2x_18 & IN2[48] | select_n2x_18 & (~ IN2[48]) | select_ne_18 & (~ IN2[49])  );
    wire logic pp_18_50;
    assign pp_18_50 = (select_e_18 & IN2[50] | select_2x_18 & IN2[49] | select_n2x_18 & (~ IN2[49]) | select_ne_18 & (~ IN2[50])  );
    wire logic pp_18_51;
    assign pp_18_51 = (select_e_18 & IN2[51] | select_2x_18 & IN2[50] | select_n2x_18 & (~ IN2[50]) | select_ne_18 & (~ IN2[51])  );
    wire logic pp_18_52;
    assign pp_18_52 = (select_e_18 & IN2[52] | select_2x_18 & IN2[51] | select_n2x_18 & (~ IN2[51]) | select_ne_18 & (~ IN2[52])  );
    wire logic pp_18_53;
    assign pp_18_53 = (select_e_18 & IN2[53] | select_2x_18 & IN2[52] | select_n2x_18 & (~ IN2[52]) | select_ne_18 & (~ IN2[53])  );
    wire logic pp_18_54;
    assign pp_18_54 = (select_e_18 & IN2[54] | select_2x_18 & IN2[53] | select_n2x_18 & (~ IN2[53]) | select_ne_18 & (~ IN2[54])  );
    wire logic pp_18_55;
    assign pp_18_55 = (select_e_18 & IN2[55] | select_2x_18 & IN2[54] | select_n2x_18 & (~ IN2[54]) | select_ne_18 & (~ IN2[55])  );
    wire logic pp_18_56;
    assign pp_18_56 = (select_e_18 & IN2[56] | select_2x_18 & IN2[55] | select_n2x_18 & (~ IN2[55]) | select_ne_18 & (~ IN2[56])  );
    wire logic pp_18_57;
    assign pp_18_57 = (select_e_18 & IN2[57] | select_2x_18 & IN2[56] | select_n2x_18 & (~ IN2[56]) | select_ne_18 & (~ IN2[57])  );
    wire logic pp_18_58;
    assign pp_18_58 = (select_e_18 & IN2[58] | select_2x_18 & IN2[57] | select_n2x_18 & (~ IN2[57]) | select_ne_18 & (~ IN2[58])  );
    wire logic pp_18_59;
    assign pp_18_59 = (select_e_18 & IN2[59] | select_2x_18 & IN2[58] | select_n2x_18 & (~ IN2[58]) | select_ne_18 & (~ IN2[59])  );
    wire logic pp_18_60;
    assign pp_18_60 = (select_e_18 & IN2[60] | select_2x_18 & IN2[59] | select_n2x_18 & (~ IN2[59]) | select_ne_18 & (~ IN2[60])  );
    wire logic pp_18_61;
    assign pp_18_61 = (select_e_18 & IN2[61] | select_2x_18 & IN2[60] | select_n2x_18 & (~ IN2[60]) | select_ne_18 & (~ IN2[61])  );
    wire logic pp_18_62;
    assign pp_18_62 = (select_e_18 & IN2[62] | select_2x_18 & IN2[61] | select_n2x_18 & (~ IN2[61]) | select_ne_18 & (~ IN2[62])  );
    wire logic pp_18_63;
    assign pp_18_63 = (select_e_18 & IN2[63] | select_2x_18 & IN2[62] | select_n2x_18 & (~ IN2[62]) | select_ne_18 & (~ IN2[63])  );
    wire logic pp_18_64;
    assign pp_18_64 = (select_e_18 & IN2[63] | select_2x_18 & IN2[63] | select_n2x_18 & (~ IN2[63]) | select_ne_18 & (~ IN2[63])  );
    wire logic pp_18_65;
    assign pp_18_65 = ~ (select_e_18 & IN2[63] | select_2x_18 & IN2[63] | select_n2x_18 & (~ IN2[63]) | select_ne_18 & (~ IN2[63])  );
    assign tcomp18 = select_ne_18 | select_n2x_18;
    
    // Signed Booth Radix-4 Partial Products Row 20
    wire logic select_e_19, select_ne_19, select_2x_19, tcomp19, select_n2x_19;
    assign select_e_19 = ((~ IN1[39]) & (IN1[38] ^ IN1[37]));
    assign select_ne_19 = IN1[39] &  (IN1[38] ^ IN1[37]);
    assign select_2x_19 = (~ IN1[39]) & IN1[38] & IN1[37];
    assign select_n2x_19 = IN1[39] & (~ IN1[38]) & (~ IN1[37]);
    wire logic pp_19_0;
    assign pp_19_0 = (select_e_19 & IN2[0] | select_2x_19 & 1'b0 | select_n2x_19 & 1'b1 | select_ne_19 & (~ IN2[0])  );
    wire logic pp_19_1;
    assign pp_19_1 = (select_e_19 & IN2[1] | select_2x_19 & IN2[0] | select_n2x_19 & (~ IN2[0]) | select_ne_19 & (~ IN2[1])  );
    wire logic pp_19_2;
    assign pp_19_2 = (select_e_19 & IN2[2] | select_2x_19 & IN2[1] | select_n2x_19 & (~ IN2[1]) | select_ne_19 & (~ IN2[2])  );
    wire logic pp_19_3;
    assign pp_19_3 = (select_e_19 & IN2[3] | select_2x_19 & IN2[2] | select_n2x_19 & (~ IN2[2]) | select_ne_19 & (~ IN2[3])  );
    wire logic pp_19_4;
    assign pp_19_4 = (select_e_19 & IN2[4] | select_2x_19 & IN2[3] | select_n2x_19 & (~ IN2[3]) | select_ne_19 & (~ IN2[4])  );
    wire logic pp_19_5;
    assign pp_19_5 = (select_e_19 & IN2[5] | select_2x_19 & IN2[4] | select_n2x_19 & (~ IN2[4]) | select_ne_19 & (~ IN2[5])  );
    wire logic pp_19_6;
    assign pp_19_6 = (select_e_19 & IN2[6] | select_2x_19 & IN2[5] | select_n2x_19 & (~ IN2[5]) | select_ne_19 & (~ IN2[6])  );
    wire logic pp_19_7;
    assign pp_19_7 = (select_e_19 & IN2[7] | select_2x_19 & IN2[6] | select_n2x_19 & (~ IN2[6]) | select_ne_19 & (~ IN2[7])  );
    wire logic pp_19_8;
    assign pp_19_8 = (select_e_19 & IN2[8] | select_2x_19 & IN2[7] | select_n2x_19 & (~ IN2[7]) | select_ne_19 & (~ IN2[8])  );
    wire logic pp_19_9;
    assign pp_19_9 = (select_e_19 & IN2[9] | select_2x_19 & IN2[8] | select_n2x_19 & (~ IN2[8]) | select_ne_19 & (~ IN2[9])  );
    wire logic pp_19_10;
    assign pp_19_10 = (select_e_19 & IN2[10] | select_2x_19 & IN2[9] | select_n2x_19 & (~ IN2[9]) | select_ne_19 & (~ IN2[10])  );
    wire logic pp_19_11;
    assign pp_19_11 = (select_e_19 & IN2[11] | select_2x_19 & IN2[10] | select_n2x_19 & (~ IN2[10]) | select_ne_19 & (~ IN2[11])  );
    wire logic pp_19_12;
    assign pp_19_12 = (select_e_19 & IN2[12] | select_2x_19 & IN2[11] | select_n2x_19 & (~ IN2[11]) | select_ne_19 & (~ IN2[12])  );
    wire logic pp_19_13;
    assign pp_19_13 = (select_e_19 & IN2[13] | select_2x_19 & IN2[12] | select_n2x_19 & (~ IN2[12]) | select_ne_19 & (~ IN2[13])  );
    wire logic pp_19_14;
    assign pp_19_14 = (select_e_19 & IN2[14] | select_2x_19 & IN2[13] | select_n2x_19 & (~ IN2[13]) | select_ne_19 & (~ IN2[14])  );
    wire logic pp_19_15;
    assign pp_19_15 = (select_e_19 & IN2[15] | select_2x_19 & IN2[14] | select_n2x_19 & (~ IN2[14]) | select_ne_19 & (~ IN2[15])  );
    wire logic pp_19_16;
    assign pp_19_16 = (select_e_19 & IN2[16] | select_2x_19 & IN2[15] | select_n2x_19 & (~ IN2[15]) | select_ne_19 & (~ IN2[16])  );
    wire logic pp_19_17;
    assign pp_19_17 = (select_e_19 & IN2[17] | select_2x_19 & IN2[16] | select_n2x_19 & (~ IN2[16]) | select_ne_19 & (~ IN2[17])  );
    wire logic pp_19_18;
    assign pp_19_18 = (select_e_19 & IN2[18] | select_2x_19 & IN2[17] | select_n2x_19 & (~ IN2[17]) | select_ne_19 & (~ IN2[18])  );
    wire logic pp_19_19;
    assign pp_19_19 = (select_e_19 & IN2[19] | select_2x_19 & IN2[18] | select_n2x_19 & (~ IN2[18]) | select_ne_19 & (~ IN2[19])  );
    wire logic pp_19_20;
    assign pp_19_20 = (select_e_19 & IN2[20] | select_2x_19 & IN2[19] | select_n2x_19 & (~ IN2[19]) | select_ne_19 & (~ IN2[20])  );
    wire logic pp_19_21;
    assign pp_19_21 = (select_e_19 & IN2[21] | select_2x_19 & IN2[20] | select_n2x_19 & (~ IN2[20]) | select_ne_19 & (~ IN2[21])  );
    wire logic pp_19_22;
    assign pp_19_22 = (select_e_19 & IN2[22] | select_2x_19 & IN2[21] | select_n2x_19 & (~ IN2[21]) | select_ne_19 & (~ IN2[22])  );
    wire logic pp_19_23;
    assign pp_19_23 = (select_e_19 & IN2[23] | select_2x_19 & IN2[22] | select_n2x_19 & (~ IN2[22]) | select_ne_19 & (~ IN2[23])  );
    wire logic pp_19_24;
    assign pp_19_24 = (select_e_19 & IN2[24] | select_2x_19 & IN2[23] | select_n2x_19 & (~ IN2[23]) | select_ne_19 & (~ IN2[24])  );
    wire logic pp_19_25;
    assign pp_19_25 = (select_e_19 & IN2[25] | select_2x_19 & IN2[24] | select_n2x_19 & (~ IN2[24]) | select_ne_19 & (~ IN2[25])  );
    wire logic pp_19_26;
    assign pp_19_26 = (select_e_19 & IN2[26] | select_2x_19 & IN2[25] | select_n2x_19 & (~ IN2[25]) | select_ne_19 & (~ IN2[26])  );
    wire logic pp_19_27;
    assign pp_19_27 = (select_e_19 & IN2[27] | select_2x_19 & IN2[26] | select_n2x_19 & (~ IN2[26]) | select_ne_19 & (~ IN2[27])  );
    wire logic pp_19_28;
    assign pp_19_28 = (select_e_19 & IN2[28] | select_2x_19 & IN2[27] | select_n2x_19 & (~ IN2[27]) | select_ne_19 & (~ IN2[28])  );
    wire logic pp_19_29;
    assign pp_19_29 = (select_e_19 & IN2[29] | select_2x_19 & IN2[28] | select_n2x_19 & (~ IN2[28]) | select_ne_19 & (~ IN2[29])  );
    wire logic pp_19_30;
    assign pp_19_30 = (select_e_19 & IN2[30] | select_2x_19 & IN2[29] | select_n2x_19 & (~ IN2[29]) | select_ne_19 & (~ IN2[30])  );
    wire logic pp_19_31;
    assign pp_19_31 = (select_e_19 & IN2[31] | select_2x_19 & IN2[30] | select_n2x_19 & (~ IN2[30]) | select_ne_19 & (~ IN2[31])  );
    wire logic pp_19_32;
    assign pp_19_32 = (select_e_19 & IN2[32] | select_2x_19 & IN2[31] | select_n2x_19 & (~ IN2[31]) | select_ne_19 & (~ IN2[32])  );
    wire logic pp_19_33;
    assign pp_19_33 = (select_e_19 & IN2[33] | select_2x_19 & IN2[32] | select_n2x_19 & (~ IN2[32]) | select_ne_19 & (~ IN2[33])  );
    wire logic pp_19_34;
    assign pp_19_34 = (select_e_19 & IN2[34] | select_2x_19 & IN2[33] | select_n2x_19 & (~ IN2[33]) | select_ne_19 & (~ IN2[34])  );
    wire logic pp_19_35;
    assign pp_19_35 = (select_e_19 & IN2[35] | select_2x_19 & IN2[34] | select_n2x_19 & (~ IN2[34]) | select_ne_19 & (~ IN2[35])  );
    wire logic pp_19_36;
    assign pp_19_36 = (select_e_19 & IN2[36] | select_2x_19 & IN2[35] | select_n2x_19 & (~ IN2[35]) | select_ne_19 & (~ IN2[36])  );
    wire logic pp_19_37;
    assign pp_19_37 = (select_e_19 & IN2[37] | select_2x_19 & IN2[36] | select_n2x_19 & (~ IN2[36]) | select_ne_19 & (~ IN2[37])  );
    wire logic pp_19_38;
    assign pp_19_38 = (select_e_19 & IN2[38] | select_2x_19 & IN2[37] | select_n2x_19 & (~ IN2[37]) | select_ne_19 & (~ IN2[38])  );
    wire logic pp_19_39;
    assign pp_19_39 = (select_e_19 & IN2[39] | select_2x_19 & IN2[38] | select_n2x_19 & (~ IN2[38]) | select_ne_19 & (~ IN2[39])  );
    wire logic pp_19_40;
    assign pp_19_40 = (select_e_19 & IN2[40] | select_2x_19 & IN2[39] | select_n2x_19 & (~ IN2[39]) | select_ne_19 & (~ IN2[40])  );
    wire logic pp_19_41;
    assign pp_19_41 = (select_e_19 & IN2[41] | select_2x_19 & IN2[40] | select_n2x_19 & (~ IN2[40]) | select_ne_19 & (~ IN2[41])  );
    wire logic pp_19_42;
    assign pp_19_42 = (select_e_19 & IN2[42] | select_2x_19 & IN2[41] | select_n2x_19 & (~ IN2[41]) | select_ne_19 & (~ IN2[42])  );
    wire logic pp_19_43;
    assign pp_19_43 = (select_e_19 & IN2[43] | select_2x_19 & IN2[42] | select_n2x_19 & (~ IN2[42]) | select_ne_19 & (~ IN2[43])  );
    wire logic pp_19_44;
    assign pp_19_44 = (select_e_19 & IN2[44] | select_2x_19 & IN2[43] | select_n2x_19 & (~ IN2[43]) | select_ne_19 & (~ IN2[44])  );
    wire logic pp_19_45;
    assign pp_19_45 = (select_e_19 & IN2[45] | select_2x_19 & IN2[44] | select_n2x_19 & (~ IN2[44]) | select_ne_19 & (~ IN2[45])  );
    wire logic pp_19_46;
    assign pp_19_46 = (select_e_19 & IN2[46] | select_2x_19 & IN2[45] | select_n2x_19 & (~ IN2[45]) | select_ne_19 & (~ IN2[46])  );
    wire logic pp_19_47;
    assign pp_19_47 = (select_e_19 & IN2[47] | select_2x_19 & IN2[46] | select_n2x_19 & (~ IN2[46]) | select_ne_19 & (~ IN2[47])  );
    wire logic pp_19_48;
    assign pp_19_48 = (select_e_19 & IN2[48] | select_2x_19 & IN2[47] | select_n2x_19 & (~ IN2[47]) | select_ne_19 & (~ IN2[48])  );
    wire logic pp_19_49;
    assign pp_19_49 = (select_e_19 & IN2[49] | select_2x_19 & IN2[48] | select_n2x_19 & (~ IN2[48]) | select_ne_19 & (~ IN2[49])  );
    wire logic pp_19_50;
    assign pp_19_50 = (select_e_19 & IN2[50] | select_2x_19 & IN2[49] | select_n2x_19 & (~ IN2[49]) | select_ne_19 & (~ IN2[50])  );
    wire logic pp_19_51;
    assign pp_19_51 = (select_e_19 & IN2[51] | select_2x_19 & IN2[50] | select_n2x_19 & (~ IN2[50]) | select_ne_19 & (~ IN2[51])  );
    wire logic pp_19_52;
    assign pp_19_52 = (select_e_19 & IN2[52] | select_2x_19 & IN2[51] | select_n2x_19 & (~ IN2[51]) | select_ne_19 & (~ IN2[52])  );
    wire logic pp_19_53;
    assign pp_19_53 = (select_e_19 & IN2[53] | select_2x_19 & IN2[52] | select_n2x_19 & (~ IN2[52]) | select_ne_19 & (~ IN2[53])  );
    wire logic pp_19_54;
    assign pp_19_54 = (select_e_19 & IN2[54] | select_2x_19 & IN2[53] | select_n2x_19 & (~ IN2[53]) | select_ne_19 & (~ IN2[54])  );
    wire logic pp_19_55;
    assign pp_19_55 = (select_e_19 & IN2[55] | select_2x_19 & IN2[54] | select_n2x_19 & (~ IN2[54]) | select_ne_19 & (~ IN2[55])  );
    wire logic pp_19_56;
    assign pp_19_56 = (select_e_19 & IN2[56] | select_2x_19 & IN2[55] | select_n2x_19 & (~ IN2[55]) | select_ne_19 & (~ IN2[56])  );
    wire logic pp_19_57;
    assign pp_19_57 = (select_e_19 & IN2[57] | select_2x_19 & IN2[56] | select_n2x_19 & (~ IN2[56]) | select_ne_19 & (~ IN2[57])  );
    wire logic pp_19_58;
    assign pp_19_58 = (select_e_19 & IN2[58] | select_2x_19 & IN2[57] | select_n2x_19 & (~ IN2[57]) | select_ne_19 & (~ IN2[58])  );
    wire logic pp_19_59;
    assign pp_19_59 = (select_e_19 & IN2[59] | select_2x_19 & IN2[58] | select_n2x_19 & (~ IN2[58]) | select_ne_19 & (~ IN2[59])  );
    wire logic pp_19_60;
    assign pp_19_60 = (select_e_19 & IN2[60] | select_2x_19 & IN2[59] | select_n2x_19 & (~ IN2[59]) | select_ne_19 & (~ IN2[60])  );
    wire logic pp_19_61;
    assign pp_19_61 = (select_e_19 & IN2[61] | select_2x_19 & IN2[60] | select_n2x_19 & (~ IN2[60]) | select_ne_19 & (~ IN2[61])  );
    wire logic pp_19_62;
    assign pp_19_62 = (select_e_19 & IN2[62] | select_2x_19 & IN2[61] | select_n2x_19 & (~ IN2[61]) | select_ne_19 & (~ IN2[62])  );
    wire logic pp_19_63;
    assign pp_19_63 = (select_e_19 & IN2[63] | select_2x_19 & IN2[62] | select_n2x_19 & (~ IN2[62]) | select_ne_19 & (~ IN2[63])  );
    wire logic pp_19_64;
    assign pp_19_64 = (select_e_19 & IN2[63] | select_2x_19 & IN2[63] | select_n2x_19 & (~ IN2[63]) | select_ne_19 & (~ IN2[63])  );
    wire logic pp_19_65;
    assign pp_19_65 = ~ (select_e_19 & IN2[63] | select_2x_19 & IN2[63] | select_n2x_19 & (~ IN2[63]) | select_ne_19 & (~ IN2[63])  );
    assign tcomp19 = select_ne_19 | select_n2x_19;
    
    // Signed Booth Radix-4 Partial Products Row 21
    wire logic select_e_20, select_ne_20, select_2x_20, tcomp20, select_n2x_20;
    assign select_e_20 = ((~ IN1[41]) & (IN1[40] ^ IN1[39]));
    assign select_ne_20 = IN1[41] &  (IN1[40] ^ IN1[39]);
    assign select_2x_20 = (~ IN1[41]) & IN1[40] & IN1[39];
    assign select_n2x_20 = IN1[41] & (~ IN1[40]) & (~ IN1[39]);
    wire logic pp_20_0;
    assign pp_20_0 = (select_e_20 & IN2[0] | select_2x_20 & 1'b0 | select_n2x_20 & 1'b1 | select_ne_20 & (~ IN2[0])  );
    wire logic pp_20_1;
    assign pp_20_1 = (select_e_20 & IN2[1] | select_2x_20 & IN2[0] | select_n2x_20 & (~ IN2[0]) | select_ne_20 & (~ IN2[1])  );
    wire logic pp_20_2;
    assign pp_20_2 = (select_e_20 & IN2[2] | select_2x_20 & IN2[1] | select_n2x_20 & (~ IN2[1]) | select_ne_20 & (~ IN2[2])  );
    wire logic pp_20_3;
    assign pp_20_3 = (select_e_20 & IN2[3] | select_2x_20 & IN2[2] | select_n2x_20 & (~ IN2[2]) | select_ne_20 & (~ IN2[3])  );
    wire logic pp_20_4;
    assign pp_20_4 = (select_e_20 & IN2[4] | select_2x_20 & IN2[3] | select_n2x_20 & (~ IN2[3]) | select_ne_20 & (~ IN2[4])  );
    wire logic pp_20_5;
    assign pp_20_5 = (select_e_20 & IN2[5] | select_2x_20 & IN2[4] | select_n2x_20 & (~ IN2[4]) | select_ne_20 & (~ IN2[5])  );
    wire logic pp_20_6;
    assign pp_20_6 = (select_e_20 & IN2[6] | select_2x_20 & IN2[5] | select_n2x_20 & (~ IN2[5]) | select_ne_20 & (~ IN2[6])  );
    wire logic pp_20_7;
    assign pp_20_7 = (select_e_20 & IN2[7] | select_2x_20 & IN2[6] | select_n2x_20 & (~ IN2[6]) | select_ne_20 & (~ IN2[7])  );
    wire logic pp_20_8;
    assign pp_20_8 = (select_e_20 & IN2[8] | select_2x_20 & IN2[7] | select_n2x_20 & (~ IN2[7]) | select_ne_20 & (~ IN2[8])  );
    wire logic pp_20_9;
    assign pp_20_9 = (select_e_20 & IN2[9] | select_2x_20 & IN2[8] | select_n2x_20 & (~ IN2[8]) | select_ne_20 & (~ IN2[9])  );
    wire logic pp_20_10;
    assign pp_20_10 = (select_e_20 & IN2[10] | select_2x_20 & IN2[9] | select_n2x_20 & (~ IN2[9]) | select_ne_20 & (~ IN2[10])  );
    wire logic pp_20_11;
    assign pp_20_11 = (select_e_20 & IN2[11] | select_2x_20 & IN2[10] | select_n2x_20 & (~ IN2[10]) | select_ne_20 & (~ IN2[11])  );
    wire logic pp_20_12;
    assign pp_20_12 = (select_e_20 & IN2[12] | select_2x_20 & IN2[11] | select_n2x_20 & (~ IN2[11]) | select_ne_20 & (~ IN2[12])  );
    wire logic pp_20_13;
    assign pp_20_13 = (select_e_20 & IN2[13] | select_2x_20 & IN2[12] | select_n2x_20 & (~ IN2[12]) | select_ne_20 & (~ IN2[13])  );
    wire logic pp_20_14;
    assign pp_20_14 = (select_e_20 & IN2[14] | select_2x_20 & IN2[13] | select_n2x_20 & (~ IN2[13]) | select_ne_20 & (~ IN2[14])  );
    wire logic pp_20_15;
    assign pp_20_15 = (select_e_20 & IN2[15] | select_2x_20 & IN2[14] | select_n2x_20 & (~ IN2[14]) | select_ne_20 & (~ IN2[15])  );
    wire logic pp_20_16;
    assign pp_20_16 = (select_e_20 & IN2[16] | select_2x_20 & IN2[15] | select_n2x_20 & (~ IN2[15]) | select_ne_20 & (~ IN2[16])  );
    wire logic pp_20_17;
    assign pp_20_17 = (select_e_20 & IN2[17] | select_2x_20 & IN2[16] | select_n2x_20 & (~ IN2[16]) | select_ne_20 & (~ IN2[17])  );
    wire logic pp_20_18;
    assign pp_20_18 = (select_e_20 & IN2[18] | select_2x_20 & IN2[17] | select_n2x_20 & (~ IN2[17]) | select_ne_20 & (~ IN2[18])  );
    wire logic pp_20_19;
    assign pp_20_19 = (select_e_20 & IN2[19] | select_2x_20 & IN2[18] | select_n2x_20 & (~ IN2[18]) | select_ne_20 & (~ IN2[19])  );
    wire logic pp_20_20;
    assign pp_20_20 = (select_e_20 & IN2[20] | select_2x_20 & IN2[19] | select_n2x_20 & (~ IN2[19]) | select_ne_20 & (~ IN2[20])  );
    wire logic pp_20_21;
    assign pp_20_21 = (select_e_20 & IN2[21] | select_2x_20 & IN2[20] | select_n2x_20 & (~ IN2[20]) | select_ne_20 & (~ IN2[21])  );
    wire logic pp_20_22;
    assign pp_20_22 = (select_e_20 & IN2[22] | select_2x_20 & IN2[21] | select_n2x_20 & (~ IN2[21]) | select_ne_20 & (~ IN2[22])  );
    wire logic pp_20_23;
    assign pp_20_23 = (select_e_20 & IN2[23] | select_2x_20 & IN2[22] | select_n2x_20 & (~ IN2[22]) | select_ne_20 & (~ IN2[23])  );
    wire logic pp_20_24;
    assign pp_20_24 = (select_e_20 & IN2[24] | select_2x_20 & IN2[23] | select_n2x_20 & (~ IN2[23]) | select_ne_20 & (~ IN2[24])  );
    wire logic pp_20_25;
    assign pp_20_25 = (select_e_20 & IN2[25] | select_2x_20 & IN2[24] | select_n2x_20 & (~ IN2[24]) | select_ne_20 & (~ IN2[25])  );
    wire logic pp_20_26;
    assign pp_20_26 = (select_e_20 & IN2[26] | select_2x_20 & IN2[25] | select_n2x_20 & (~ IN2[25]) | select_ne_20 & (~ IN2[26])  );
    wire logic pp_20_27;
    assign pp_20_27 = (select_e_20 & IN2[27] | select_2x_20 & IN2[26] | select_n2x_20 & (~ IN2[26]) | select_ne_20 & (~ IN2[27])  );
    wire logic pp_20_28;
    assign pp_20_28 = (select_e_20 & IN2[28] | select_2x_20 & IN2[27] | select_n2x_20 & (~ IN2[27]) | select_ne_20 & (~ IN2[28])  );
    wire logic pp_20_29;
    assign pp_20_29 = (select_e_20 & IN2[29] | select_2x_20 & IN2[28] | select_n2x_20 & (~ IN2[28]) | select_ne_20 & (~ IN2[29])  );
    wire logic pp_20_30;
    assign pp_20_30 = (select_e_20 & IN2[30] | select_2x_20 & IN2[29] | select_n2x_20 & (~ IN2[29]) | select_ne_20 & (~ IN2[30])  );
    wire logic pp_20_31;
    assign pp_20_31 = (select_e_20 & IN2[31] | select_2x_20 & IN2[30] | select_n2x_20 & (~ IN2[30]) | select_ne_20 & (~ IN2[31])  );
    wire logic pp_20_32;
    assign pp_20_32 = (select_e_20 & IN2[32] | select_2x_20 & IN2[31] | select_n2x_20 & (~ IN2[31]) | select_ne_20 & (~ IN2[32])  );
    wire logic pp_20_33;
    assign pp_20_33 = (select_e_20 & IN2[33] | select_2x_20 & IN2[32] | select_n2x_20 & (~ IN2[32]) | select_ne_20 & (~ IN2[33])  );
    wire logic pp_20_34;
    assign pp_20_34 = (select_e_20 & IN2[34] | select_2x_20 & IN2[33] | select_n2x_20 & (~ IN2[33]) | select_ne_20 & (~ IN2[34])  );
    wire logic pp_20_35;
    assign pp_20_35 = (select_e_20 & IN2[35] | select_2x_20 & IN2[34] | select_n2x_20 & (~ IN2[34]) | select_ne_20 & (~ IN2[35])  );
    wire logic pp_20_36;
    assign pp_20_36 = (select_e_20 & IN2[36] | select_2x_20 & IN2[35] | select_n2x_20 & (~ IN2[35]) | select_ne_20 & (~ IN2[36])  );
    wire logic pp_20_37;
    assign pp_20_37 = (select_e_20 & IN2[37] | select_2x_20 & IN2[36] | select_n2x_20 & (~ IN2[36]) | select_ne_20 & (~ IN2[37])  );
    wire logic pp_20_38;
    assign pp_20_38 = (select_e_20 & IN2[38] | select_2x_20 & IN2[37] | select_n2x_20 & (~ IN2[37]) | select_ne_20 & (~ IN2[38])  );
    wire logic pp_20_39;
    assign pp_20_39 = (select_e_20 & IN2[39] | select_2x_20 & IN2[38] | select_n2x_20 & (~ IN2[38]) | select_ne_20 & (~ IN2[39])  );
    wire logic pp_20_40;
    assign pp_20_40 = (select_e_20 & IN2[40] | select_2x_20 & IN2[39] | select_n2x_20 & (~ IN2[39]) | select_ne_20 & (~ IN2[40])  );
    wire logic pp_20_41;
    assign pp_20_41 = (select_e_20 & IN2[41] | select_2x_20 & IN2[40] | select_n2x_20 & (~ IN2[40]) | select_ne_20 & (~ IN2[41])  );
    wire logic pp_20_42;
    assign pp_20_42 = (select_e_20 & IN2[42] | select_2x_20 & IN2[41] | select_n2x_20 & (~ IN2[41]) | select_ne_20 & (~ IN2[42])  );
    wire logic pp_20_43;
    assign pp_20_43 = (select_e_20 & IN2[43] | select_2x_20 & IN2[42] | select_n2x_20 & (~ IN2[42]) | select_ne_20 & (~ IN2[43])  );
    wire logic pp_20_44;
    assign pp_20_44 = (select_e_20 & IN2[44] | select_2x_20 & IN2[43] | select_n2x_20 & (~ IN2[43]) | select_ne_20 & (~ IN2[44])  );
    wire logic pp_20_45;
    assign pp_20_45 = (select_e_20 & IN2[45] | select_2x_20 & IN2[44] | select_n2x_20 & (~ IN2[44]) | select_ne_20 & (~ IN2[45])  );
    wire logic pp_20_46;
    assign pp_20_46 = (select_e_20 & IN2[46] | select_2x_20 & IN2[45] | select_n2x_20 & (~ IN2[45]) | select_ne_20 & (~ IN2[46])  );
    wire logic pp_20_47;
    assign pp_20_47 = (select_e_20 & IN2[47] | select_2x_20 & IN2[46] | select_n2x_20 & (~ IN2[46]) | select_ne_20 & (~ IN2[47])  );
    wire logic pp_20_48;
    assign pp_20_48 = (select_e_20 & IN2[48] | select_2x_20 & IN2[47] | select_n2x_20 & (~ IN2[47]) | select_ne_20 & (~ IN2[48])  );
    wire logic pp_20_49;
    assign pp_20_49 = (select_e_20 & IN2[49] | select_2x_20 & IN2[48] | select_n2x_20 & (~ IN2[48]) | select_ne_20 & (~ IN2[49])  );
    wire logic pp_20_50;
    assign pp_20_50 = (select_e_20 & IN2[50] | select_2x_20 & IN2[49] | select_n2x_20 & (~ IN2[49]) | select_ne_20 & (~ IN2[50])  );
    wire logic pp_20_51;
    assign pp_20_51 = (select_e_20 & IN2[51] | select_2x_20 & IN2[50] | select_n2x_20 & (~ IN2[50]) | select_ne_20 & (~ IN2[51])  );
    wire logic pp_20_52;
    assign pp_20_52 = (select_e_20 & IN2[52] | select_2x_20 & IN2[51] | select_n2x_20 & (~ IN2[51]) | select_ne_20 & (~ IN2[52])  );
    wire logic pp_20_53;
    assign pp_20_53 = (select_e_20 & IN2[53] | select_2x_20 & IN2[52] | select_n2x_20 & (~ IN2[52]) | select_ne_20 & (~ IN2[53])  );
    wire logic pp_20_54;
    assign pp_20_54 = (select_e_20 & IN2[54] | select_2x_20 & IN2[53] | select_n2x_20 & (~ IN2[53]) | select_ne_20 & (~ IN2[54])  );
    wire logic pp_20_55;
    assign pp_20_55 = (select_e_20 & IN2[55] | select_2x_20 & IN2[54] | select_n2x_20 & (~ IN2[54]) | select_ne_20 & (~ IN2[55])  );
    wire logic pp_20_56;
    assign pp_20_56 = (select_e_20 & IN2[56] | select_2x_20 & IN2[55] | select_n2x_20 & (~ IN2[55]) | select_ne_20 & (~ IN2[56])  );
    wire logic pp_20_57;
    assign pp_20_57 = (select_e_20 & IN2[57] | select_2x_20 & IN2[56] | select_n2x_20 & (~ IN2[56]) | select_ne_20 & (~ IN2[57])  );
    wire logic pp_20_58;
    assign pp_20_58 = (select_e_20 & IN2[58] | select_2x_20 & IN2[57] | select_n2x_20 & (~ IN2[57]) | select_ne_20 & (~ IN2[58])  );
    wire logic pp_20_59;
    assign pp_20_59 = (select_e_20 & IN2[59] | select_2x_20 & IN2[58] | select_n2x_20 & (~ IN2[58]) | select_ne_20 & (~ IN2[59])  );
    wire logic pp_20_60;
    assign pp_20_60 = (select_e_20 & IN2[60] | select_2x_20 & IN2[59] | select_n2x_20 & (~ IN2[59]) | select_ne_20 & (~ IN2[60])  );
    wire logic pp_20_61;
    assign pp_20_61 = (select_e_20 & IN2[61] | select_2x_20 & IN2[60] | select_n2x_20 & (~ IN2[60]) | select_ne_20 & (~ IN2[61])  );
    wire logic pp_20_62;
    assign pp_20_62 = (select_e_20 & IN2[62] | select_2x_20 & IN2[61] | select_n2x_20 & (~ IN2[61]) | select_ne_20 & (~ IN2[62])  );
    wire logic pp_20_63;
    assign pp_20_63 = (select_e_20 & IN2[63] | select_2x_20 & IN2[62] | select_n2x_20 & (~ IN2[62]) | select_ne_20 & (~ IN2[63])  );
    wire logic pp_20_64;
    assign pp_20_64 = (select_e_20 & IN2[63] | select_2x_20 & IN2[63] | select_n2x_20 & (~ IN2[63]) | select_ne_20 & (~ IN2[63])  );
    wire logic pp_20_65;
    assign pp_20_65 = ~ (select_e_20 & IN2[63] | select_2x_20 & IN2[63] | select_n2x_20 & (~ IN2[63]) | select_ne_20 & (~ IN2[63])  );
    assign tcomp20 = select_ne_20 | select_n2x_20;
    
    // Signed Booth Radix-4 Partial Products Row 22
    wire logic select_e_21, select_ne_21, select_2x_21, tcomp21, select_n2x_21;
    assign select_e_21 = ((~ IN1[43]) & (IN1[42] ^ IN1[41]));
    assign select_ne_21 = IN1[43] &  (IN1[42] ^ IN1[41]);
    assign select_2x_21 = (~ IN1[43]) & IN1[42] & IN1[41];
    assign select_n2x_21 = IN1[43] & (~ IN1[42]) & (~ IN1[41]);
    wire logic pp_21_0;
    assign pp_21_0 = (select_e_21 & IN2[0] | select_2x_21 & 1'b0 | select_n2x_21 & 1'b1 | select_ne_21 & (~ IN2[0])  );
    wire logic pp_21_1;
    assign pp_21_1 = (select_e_21 & IN2[1] | select_2x_21 & IN2[0] | select_n2x_21 & (~ IN2[0]) | select_ne_21 & (~ IN2[1])  );
    wire logic pp_21_2;
    assign pp_21_2 = (select_e_21 & IN2[2] | select_2x_21 & IN2[1] | select_n2x_21 & (~ IN2[1]) | select_ne_21 & (~ IN2[2])  );
    wire logic pp_21_3;
    assign pp_21_3 = (select_e_21 & IN2[3] | select_2x_21 & IN2[2] | select_n2x_21 & (~ IN2[2]) | select_ne_21 & (~ IN2[3])  );
    wire logic pp_21_4;
    assign pp_21_4 = (select_e_21 & IN2[4] | select_2x_21 & IN2[3] | select_n2x_21 & (~ IN2[3]) | select_ne_21 & (~ IN2[4])  );
    wire logic pp_21_5;
    assign pp_21_5 = (select_e_21 & IN2[5] | select_2x_21 & IN2[4] | select_n2x_21 & (~ IN2[4]) | select_ne_21 & (~ IN2[5])  );
    wire logic pp_21_6;
    assign pp_21_6 = (select_e_21 & IN2[6] | select_2x_21 & IN2[5] | select_n2x_21 & (~ IN2[5]) | select_ne_21 & (~ IN2[6])  );
    wire logic pp_21_7;
    assign pp_21_7 = (select_e_21 & IN2[7] | select_2x_21 & IN2[6] | select_n2x_21 & (~ IN2[6]) | select_ne_21 & (~ IN2[7])  );
    wire logic pp_21_8;
    assign pp_21_8 = (select_e_21 & IN2[8] | select_2x_21 & IN2[7] | select_n2x_21 & (~ IN2[7]) | select_ne_21 & (~ IN2[8])  );
    wire logic pp_21_9;
    assign pp_21_9 = (select_e_21 & IN2[9] | select_2x_21 & IN2[8] | select_n2x_21 & (~ IN2[8]) | select_ne_21 & (~ IN2[9])  );
    wire logic pp_21_10;
    assign pp_21_10 = (select_e_21 & IN2[10] | select_2x_21 & IN2[9] | select_n2x_21 & (~ IN2[9]) | select_ne_21 & (~ IN2[10])  );
    wire logic pp_21_11;
    assign pp_21_11 = (select_e_21 & IN2[11] | select_2x_21 & IN2[10] | select_n2x_21 & (~ IN2[10]) | select_ne_21 & (~ IN2[11])  );
    wire logic pp_21_12;
    assign pp_21_12 = (select_e_21 & IN2[12] | select_2x_21 & IN2[11] | select_n2x_21 & (~ IN2[11]) | select_ne_21 & (~ IN2[12])  );
    wire logic pp_21_13;
    assign pp_21_13 = (select_e_21 & IN2[13] | select_2x_21 & IN2[12] | select_n2x_21 & (~ IN2[12]) | select_ne_21 & (~ IN2[13])  );
    wire logic pp_21_14;
    assign pp_21_14 = (select_e_21 & IN2[14] | select_2x_21 & IN2[13] | select_n2x_21 & (~ IN2[13]) | select_ne_21 & (~ IN2[14])  );
    wire logic pp_21_15;
    assign pp_21_15 = (select_e_21 & IN2[15] | select_2x_21 & IN2[14] | select_n2x_21 & (~ IN2[14]) | select_ne_21 & (~ IN2[15])  );
    wire logic pp_21_16;
    assign pp_21_16 = (select_e_21 & IN2[16] | select_2x_21 & IN2[15] | select_n2x_21 & (~ IN2[15]) | select_ne_21 & (~ IN2[16])  );
    wire logic pp_21_17;
    assign pp_21_17 = (select_e_21 & IN2[17] | select_2x_21 & IN2[16] | select_n2x_21 & (~ IN2[16]) | select_ne_21 & (~ IN2[17])  );
    wire logic pp_21_18;
    assign pp_21_18 = (select_e_21 & IN2[18] | select_2x_21 & IN2[17] | select_n2x_21 & (~ IN2[17]) | select_ne_21 & (~ IN2[18])  );
    wire logic pp_21_19;
    assign pp_21_19 = (select_e_21 & IN2[19] | select_2x_21 & IN2[18] | select_n2x_21 & (~ IN2[18]) | select_ne_21 & (~ IN2[19])  );
    wire logic pp_21_20;
    assign pp_21_20 = (select_e_21 & IN2[20] | select_2x_21 & IN2[19] | select_n2x_21 & (~ IN2[19]) | select_ne_21 & (~ IN2[20])  );
    wire logic pp_21_21;
    assign pp_21_21 = (select_e_21 & IN2[21] | select_2x_21 & IN2[20] | select_n2x_21 & (~ IN2[20]) | select_ne_21 & (~ IN2[21])  );
    wire logic pp_21_22;
    assign pp_21_22 = (select_e_21 & IN2[22] | select_2x_21 & IN2[21] | select_n2x_21 & (~ IN2[21]) | select_ne_21 & (~ IN2[22])  );
    wire logic pp_21_23;
    assign pp_21_23 = (select_e_21 & IN2[23] | select_2x_21 & IN2[22] | select_n2x_21 & (~ IN2[22]) | select_ne_21 & (~ IN2[23])  );
    wire logic pp_21_24;
    assign pp_21_24 = (select_e_21 & IN2[24] | select_2x_21 & IN2[23] | select_n2x_21 & (~ IN2[23]) | select_ne_21 & (~ IN2[24])  );
    wire logic pp_21_25;
    assign pp_21_25 = (select_e_21 & IN2[25] | select_2x_21 & IN2[24] | select_n2x_21 & (~ IN2[24]) | select_ne_21 & (~ IN2[25])  );
    wire logic pp_21_26;
    assign pp_21_26 = (select_e_21 & IN2[26] | select_2x_21 & IN2[25] | select_n2x_21 & (~ IN2[25]) | select_ne_21 & (~ IN2[26])  );
    wire logic pp_21_27;
    assign pp_21_27 = (select_e_21 & IN2[27] | select_2x_21 & IN2[26] | select_n2x_21 & (~ IN2[26]) | select_ne_21 & (~ IN2[27])  );
    wire logic pp_21_28;
    assign pp_21_28 = (select_e_21 & IN2[28] | select_2x_21 & IN2[27] | select_n2x_21 & (~ IN2[27]) | select_ne_21 & (~ IN2[28])  );
    wire logic pp_21_29;
    assign pp_21_29 = (select_e_21 & IN2[29] | select_2x_21 & IN2[28] | select_n2x_21 & (~ IN2[28]) | select_ne_21 & (~ IN2[29])  );
    wire logic pp_21_30;
    assign pp_21_30 = (select_e_21 & IN2[30] | select_2x_21 & IN2[29] | select_n2x_21 & (~ IN2[29]) | select_ne_21 & (~ IN2[30])  );
    wire logic pp_21_31;
    assign pp_21_31 = (select_e_21 & IN2[31] | select_2x_21 & IN2[30] | select_n2x_21 & (~ IN2[30]) | select_ne_21 & (~ IN2[31])  );
    wire logic pp_21_32;
    assign pp_21_32 = (select_e_21 & IN2[32] | select_2x_21 & IN2[31] | select_n2x_21 & (~ IN2[31]) | select_ne_21 & (~ IN2[32])  );
    wire logic pp_21_33;
    assign pp_21_33 = (select_e_21 & IN2[33] | select_2x_21 & IN2[32] | select_n2x_21 & (~ IN2[32]) | select_ne_21 & (~ IN2[33])  );
    wire logic pp_21_34;
    assign pp_21_34 = (select_e_21 & IN2[34] | select_2x_21 & IN2[33] | select_n2x_21 & (~ IN2[33]) | select_ne_21 & (~ IN2[34])  );
    wire logic pp_21_35;
    assign pp_21_35 = (select_e_21 & IN2[35] | select_2x_21 & IN2[34] | select_n2x_21 & (~ IN2[34]) | select_ne_21 & (~ IN2[35])  );
    wire logic pp_21_36;
    assign pp_21_36 = (select_e_21 & IN2[36] | select_2x_21 & IN2[35] | select_n2x_21 & (~ IN2[35]) | select_ne_21 & (~ IN2[36])  );
    wire logic pp_21_37;
    assign pp_21_37 = (select_e_21 & IN2[37] | select_2x_21 & IN2[36] | select_n2x_21 & (~ IN2[36]) | select_ne_21 & (~ IN2[37])  );
    wire logic pp_21_38;
    assign pp_21_38 = (select_e_21 & IN2[38] | select_2x_21 & IN2[37] | select_n2x_21 & (~ IN2[37]) | select_ne_21 & (~ IN2[38])  );
    wire logic pp_21_39;
    assign pp_21_39 = (select_e_21 & IN2[39] | select_2x_21 & IN2[38] | select_n2x_21 & (~ IN2[38]) | select_ne_21 & (~ IN2[39])  );
    wire logic pp_21_40;
    assign pp_21_40 = (select_e_21 & IN2[40] | select_2x_21 & IN2[39] | select_n2x_21 & (~ IN2[39]) | select_ne_21 & (~ IN2[40])  );
    wire logic pp_21_41;
    assign pp_21_41 = (select_e_21 & IN2[41] | select_2x_21 & IN2[40] | select_n2x_21 & (~ IN2[40]) | select_ne_21 & (~ IN2[41])  );
    wire logic pp_21_42;
    assign pp_21_42 = (select_e_21 & IN2[42] | select_2x_21 & IN2[41] | select_n2x_21 & (~ IN2[41]) | select_ne_21 & (~ IN2[42])  );
    wire logic pp_21_43;
    assign pp_21_43 = (select_e_21 & IN2[43] | select_2x_21 & IN2[42] | select_n2x_21 & (~ IN2[42]) | select_ne_21 & (~ IN2[43])  );
    wire logic pp_21_44;
    assign pp_21_44 = (select_e_21 & IN2[44] | select_2x_21 & IN2[43] | select_n2x_21 & (~ IN2[43]) | select_ne_21 & (~ IN2[44])  );
    wire logic pp_21_45;
    assign pp_21_45 = (select_e_21 & IN2[45] | select_2x_21 & IN2[44] | select_n2x_21 & (~ IN2[44]) | select_ne_21 & (~ IN2[45])  );
    wire logic pp_21_46;
    assign pp_21_46 = (select_e_21 & IN2[46] | select_2x_21 & IN2[45] | select_n2x_21 & (~ IN2[45]) | select_ne_21 & (~ IN2[46])  );
    wire logic pp_21_47;
    assign pp_21_47 = (select_e_21 & IN2[47] | select_2x_21 & IN2[46] | select_n2x_21 & (~ IN2[46]) | select_ne_21 & (~ IN2[47])  );
    wire logic pp_21_48;
    assign pp_21_48 = (select_e_21 & IN2[48] | select_2x_21 & IN2[47] | select_n2x_21 & (~ IN2[47]) | select_ne_21 & (~ IN2[48])  );
    wire logic pp_21_49;
    assign pp_21_49 = (select_e_21 & IN2[49] | select_2x_21 & IN2[48] | select_n2x_21 & (~ IN2[48]) | select_ne_21 & (~ IN2[49])  );
    wire logic pp_21_50;
    assign pp_21_50 = (select_e_21 & IN2[50] | select_2x_21 & IN2[49] | select_n2x_21 & (~ IN2[49]) | select_ne_21 & (~ IN2[50])  );
    wire logic pp_21_51;
    assign pp_21_51 = (select_e_21 & IN2[51] | select_2x_21 & IN2[50] | select_n2x_21 & (~ IN2[50]) | select_ne_21 & (~ IN2[51])  );
    wire logic pp_21_52;
    assign pp_21_52 = (select_e_21 & IN2[52] | select_2x_21 & IN2[51] | select_n2x_21 & (~ IN2[51]) | select_ne_21 & (~ IN2[52])  );
    wire logic pp_21_53;
    assign pp_21_53 = (select_e_21 & IN2[53] | select_2x_21 & IN2[52] | select_n2x_21 & (~ IN2[52]) | select_ne_21 & (~ IN2[53])  );
    wire logic pp_21_54;
    assign pp_21_54 = (select_e_21 & IN2[54] | select_2x_21 & IN2[53] | select_n2x_21 & (~ IN2[53]) | select_ne_21 & (~ IN2[54])  );
    wire logic pp_21_55;
    assign pp_21_55 = (select_e_21 & IN2[55] | select_2x_21 & IN2[54] | select_n2x_21 & (~ IN2[54]) | select_ne_21 & (~ IN2[55])  );
    wire logic pp_21_56;
    assign pp_21_56 = (select_e_21 & IN2[56] | select_2x_21 & IN2[55] | select_n2x_21 & (~ IN2[55]) | select_ne_21 & (~ IN2[56])  );
    wire logic pp_21_57;
    assign pp_21_57 = (select_e_21 & IN2[57] | select_2x_21 & IN2[56] | select_n2x_21 & (~ IN2[56]) | select_ne_21 & (~ IN2[57])  );
    wire logic pp_21_58;
    assign pp_21_58 = (select_e_21 & IN2[58] | select_2x_21 & IN2[57] | select_n2x_21 & (~ IN2[57]) | select_ne_21 & (~ IN2[58])  );
    wire logic pp_21_59;
    assign pp_21_59 = (select_e_21 & IN2[59] | select_2x_21 & IN2[58] | select_n2x_21 & (~ IN2[58]) | select_ne_21 & (~ IN2[59])  );
    wire logic pp_21_60;
    assign pp_21_60 = (select_e_21 & IN2[60] | select_2x_21 & IN2[59] | select_n2x_21 & (~ IN2[59]) | select_ne_21 & (~ IN2[60])  );
    wire logic pp_21_61;
    assign pp_21_61 = (select_e_21 & IN2[61] | select_2x_21 & IN2[60] | select_n2x_21 & (~ IN2[60]) | select_ne_21 & (~ IN2[61])  );
    wire logic pp_21_62;
    assign pp_21_62 = (select_e_21 & IN2[62] | select_2x_21 & IN2[61] | select_n2x_21 & (~ IN2[61]) | select_ne_21 & (~ IN2[62])  );
    wire logic pp_21_63;
    assign pp_21_63 = (select_e_21 & IN2[63] | select_2x_21 & IN2[62] | select_n2x_21 & (~ IN2[62]) | select_ne_21 & (~ IN2[63])  );
    wire logic pp_21_64;
    assign pp_21_64 = (select_e_21 & IN2[63] | select_2x_21 & IN2[63] | select_n2x_21 & (~ IN2[63]) | select_ne_21 & (~ IN2[63])  );
    wire logic pp_21_65;
    assign pp_21_65 = ~ (select_e_21 & IN2[63] | select_2x_21 & IN2[63] | select_n2x_21 & (~ IN2[63]) | select_ne_21 & (~ IN2[63])  );
    assign tcomp21 = select_ne_21 | select_n2x_21;
    
    // Signed Booth Radix-4 Partial Products Row 23
    wire logic select_e_22, select_ne_22, select_2x_22, tcomp22, select_n2x_22;
    assign select_e_22 = ((~ IN1[45]) & (IN1[44] ^ IN1[43]));
    assign select_ne_22 = IN1[45] &  (IN1[44] ^ IN1[43]);
    assign select_2x_22 = (~ IN1[45]) & IN1[44] & IN1[43];
    assign select_n2x_22 = IN1[45] & (~ IN1[44]) & (~ IN1[43]);
    wire logic pp_22_0;
    assign pp_22_0 = (select_e_22 & IN2[0] | select_2x_22 & 1'b0 | select_n2x_22 & 1'b1 | select_ne_22 & (~ IN2[0])  );
    wire logic pp_22_1;
    assign pp_22_1 = (select_e_22 & IN2[1] | select_2x_22 & IN2[0] | select_n2x_22 & (~ IN2[0]) | select_ne_22 & (~ IN2[1])  );
    wire logic pp_22_2;
    assign pp_22_2 = (select_e_22 & IN2[2] | select_2x_22 & IN2[1] | select_n2x_22 & (~ IN2[1]) | select_ne_22 & (~ IN2[2])  );
    wire logic pp_22_3;
    assign pp_22_3 = (select_e_22 & IN2[3] | select_2x_22 & IN2[2] | select_n2x_22 & (~ IN2[2]) | select_ne_22 & (~ IN2[3])  );
    wire logic pp_22_4;
    assign pp_22_4 = (select_e_22 & IN2[4] | select_2x_22 & IN2[3] | select_n2x_22 & (~ IN2[3]) | select_ne_22 & (~ IN2[4])  );
    wire logic pp_22_5;
    assign pp_22_5 = (select_e_22 & IN2[5] | select_2x_22 & IN2[4] | select_n2x_22 & (~ IN2[4]) | select_ne_22 & (~ IN2[5])  );
    wire logic pp_22_6;
    assign pp_22_6 = (select_e_22 & IN2[6] | select_2x_22 & IN2[5] | select_n2x_22 & (~ IN2[5]) | select_ne_22 & (~ IN2[6])  );
    wire logic pp_22_7;
    assign pp_22_7 = (select_e_22 & IN2[7] | select_2x_22 & IN2[6] | select_n2x_22 & (~ IN2[6]) | select_ne_22 & (~ IN2[7])  );
    wire logic pp_22_8;
    assign pp_22_8 = (select_e_22 & IN2[8] | select_2x_22 & IN2[7] | select_n2x_22 & (~ IN2[7]) | select_ne_22 & (~ IN2[8])  );
    wire logic pp_22_9;
    assign pp_22_9 = (select_e_22 & IN2[9] | select_2x_22 & IN2[8] | select_n2x_22 & (~ IN2[8]) | select_ne_22 & (~ IN2[9])  );
    wire logic pp_22_10;
    assign pp_22_10 = (select_e_22 & IN2[10] | select_2x_22 & IN2[9] | select_n2x_22 & (~ IN2[9]) | select_ne_22 & (~ IN2[10])  );
    wire logic pp_22_11;
    assign pp_22_11 = (select_e_22 & IN2[11] | select_2x_22 & IN2[10] | select_n2x_22 & (~ IN2[10]) | select_ne_22 & (~ IN2[11])  );
    wire logic pp_22_12;
    assign pp_22_12 = (select_e_22 & IN2[12] | select_2x_22 & IN2[11] | select_n2x_22 & (~ IN2[11]) | select_ne_22 & (~ IN2[12])  );
    wire logic pp_22_13;
    assign pp_22_13 = (select_e_22 & IN2[13] | select_2x_22 & IN2[12] | select_n2x_22 & (~ IN2[12]) | select_ne_22 & (~ IN2[13])  );
    wire logic pp_22_14;
    assign pp_22_14 = (select_e_22 & IN2[14] | select_2x_22 & IN2[13] | select_n2x_22 & (~ IN2[13]) | select_ne_22 & (~ IN2[14])  );
    wire logic pp_22_15;
    assign pp_22_15 = (select_e_22 & IN2[15] | select_2x_22 & IN2[14] | select_n2x_22 & (~ IN2[14]) | select_ne_22 & (~ IN2[15])  );
    wire logic pp_22_16;
    assign pp_22_16 = (select_e_22 & IN2[16] | select_2x_22 & IN2[15] | select_n2x_22 & (~ IN2[15]) | select_ne_22 & (~ IN2[16])  );
    wire logic pp_22_17;
    assign pp_22_17 = (select_e_22 & IN2[17] | select_2x_22 & IN2[16] | select_n2x_22 & (~ IN2[16]) | select_ne_22 & (~ IN2[17])  );
    wire logic pp_22_18;
    assign pp_22_18 = (select_e_22 & IN2[18] | select_2x_22 & IN2[17] | select_n2x_22 & (~ IN2[17]) | select_ne_22 & (~ IN2[18])  );
    wire logic pp_22_19;
    assign pp_22_19 = (select_e_22 & IN2[19] | select_2x_22 & IN2[18] | select_n2x_22 & (~ IN2[18]) | select_ne_22 & (~ IN2[19])  );
    wire logic pp_22_20;
    assign pp_22_20 = (select_e_22 & IN2[20] | select_2x_22 & IN2[19] | select_n2x_22 & (~ IN2[19]) | select_ne_22 & (~ IN2[20])  );
    wire logic pp_22_21;
    assign pp_22_21 = (select_e_22 & IN2[21] | select_2x_22 & IN2[20] | select_n2x_22 & (~ IN2[20]) | select_ne_22 & (~ IN2[21])  );
    wire logic pp_22_22;
    assign pp_22_22 = (select_e_22 & IN2[22] | select_2x_22 & IN2[21] | select_n2x_22 & (~ IN2[21]) | select_ne_22 & (~ IN2[22])  );
    wire logic pp_22_23;
    assign pp_22_23 = (select_e_22 & IN2[23] | select_2x_22 & IN2[22] | select_n2x_22 & (~ IN2[22]) | select_ne_22 & (~ IN2[23])  );
    wire logic pp_22_24;
    assign pp_22_24 = (select_e_22 & IN2[24] | select_2x_22 & IN2[23] | select_n2x_22 & (~ IN2[23]) | select_ne_22 & (~ IN2[24])  );
    wire logic pp_22_25;
    assign pp_22_25 = (select_e_22 & IN2[25] | select_2x_22 & IN2[24] | select_n2x_22 & (~ IN2[24]) | select_ne_22 & (~ IN2[25])  );
    wire logic pp_22_26;
    assign pp_22_26 = (select_e_22 & IN2[26] | select_2x_22 & IN2[25] | select_n2x_22 & (~ IN2[25]) | select_ne_22 & (~ IN2[26])  );
    wire logic pp_22_27;
    assign pp_22_27 = (select_e_22 & IN2[27] | select_2x_22 & IN2[26] | select_n2x_22 & (~ IN2[26]) | select_ne_22 & (~ IN2[27])  );
    wire logic pp_22_28;
    assign pp_22_28 = (select_e_22 & IN2[28] | select_2x_22 & IN2[27] | select_n2x_22 & (~ IN2[27]) | select_ne_22 & (~ IN2[28])  );
    wire logic pp_22_29;
    assign pp_22_29 = (select_e_22 & IN2[29] | select_2x_22 & IN2[28] | select_n2x_22 & (~ IN2[28]) | select_ne_22 & (~ IN2[29])  );
    wire logic pp_22_30;
    assign pp_22_30 = (select_e_22 & IN2[30] | select_2x_22 & IN2[29] | select_n2x_22 & (~ IN2[29]) | select_ne_22 & (~ IN2[30])  );
    wire logic pp_22_31;
    assign pp_22_31 = (select_e_22 & IN2[31] | select_2x_22 & IN2[30] | select_n2x_22 & (~ IN2[30]) | select_ne_22 & (~ IN2[31])  );
    wire logic pp_22_32;
    assign pp_22_32 = (select_e_22 & IN2[32] | select_2x_22 & IN2[31] | select_n2x_22 & (~ IN2[31]) | select_ne_22 & (~ IN2[32])  );
    wire logic pp_22_33;
    assign pp_22_33 = (select_e_22 & IN2[33] | select_2x_22 & IN2[32] | select_n2x_22 & (~ IN2[32]) | select_ne_22 & (~ IN2[33])  );
    wire logic pp_22_34;
    assign pp_22_34 = (select_e_22 & IN2[34] | select_2x_22 & IN2[33] | select_n2x_22 & (~ IN2[33]) | select_ne_22 & (~ IN2[34])  );
    wire logic pp_22_35;
    assign pp_22_35 = (select_e_22 & IN2[35] | select_2x_22 & IN2[34] | select_n2x_22 & (~ IN2[34]) | select_ne_22 & (~ IN2[35])  );
    wire logic pp_22_36;
    assign pp_22_36 = (select_e_22 & IN2[36] | select_2x_22 & IN2[35] | select_n2x_22 & (~ IN2[35]) | select_ne_22 & (~ IN2[36])  );
    wire logic pp_22_37;
    assign pp_22_37 = (select_e_22 & IN2[37] | select_2x_22 & IN2[36] | select_n2x_22 & (~ IN2[36]) | select_ne_22 & (~ IN2[37])  );
    wire logic pp_22_38;
    assign pp_22_38 = (select_e_22 & IN2[38] | select_2x_22 & IN2[37] | select_n2x_22 & (~ IN2[37]) | select_ne_22 & (~ IN2[38])  );
    wire logic pp_22_39;
    assign pp_22_39 = (select_e_22 & IN2[39] | select_2x_22 & IN2[38] | select_n2x_22 & (~ IN2[38]) | select_ne_22 & (~ IN2[39])  );
    wire logic pp_22_40;
    assign pp_22_40 = (select_e_22 & IN2[40] | select_2x_22 & IN2[39] | select_n2x_22 & (~ IN2[39]) | select_ne_22 & (~ IN2[40])  );
    wire logic pp_22_41;
    assign pp_22_41 = (select_e_22 & IN2[41] | select_2x_22 & IN2[40] | select_n2x_22 & (~ IN2[40]) | select_ne_22 & (~ IN2[41])  );
    wire logic pp_22_42;
    assign pp_22_42 = (select_e_22 & IN2[42] | select_2x_22 & IN2[41] | select_n2x_22 & (~ IN2[41]) | select_ne_22 & (~ IN2[42])  );
    wire logic pp_22_43;
    assign pp_22_43 = (select_e_22 & IN2[43] | select_2x_22 & IN2[42] | select_n2x_22 & (~ IN2[42]) | select_ne_22 & (~ IN2[43])  );
    wire logic pp_22_44;
    assign pp_22_44 = (select_e_22 & IN2[44] | select_2x_22 & IN2[43] | select_n2x_22 & (~ IN2[43]) | select_ne_22 & (~ IN2[44])  );
    wire logic pp_22_45;
    assign pp_22_45 = (select_e_22 & IN2[45] | select_2x_22 & IN2[44] | select_n2x_22 & (~ IN2[44]) | select_ne_22 & (~ IN2[45])  );
    wire logic pp_22_46;
    assign pp_22_46 = (select_e_22 & IN2[46] | select_2x_22 & IN2[45] | select_n2x_22 & (~ IN2[45]) | select_ne_22 & (~ IN2[46])  );
    wire logic pp_22_47;
    assign pp_22_47 = (select_e_22 & IN2[47] | select_2x_22 & IN2[46] | select_n2x_22 & (~ IN2[46]) | select_ne_22 & (~ IN2[47])  );
    wire logic pp_22_48;
    assign pp_22_48 = (select_e_22 & IN2[48] | select_2x_22 & IN2[47] | select_n2x_22 & (~ IN2[47]) | select_ne_22 & (~ IN2[48])  );
    wire logic pp_22_49;
    assign pp_22_49 = (select_e_22 & IN2[49] | select_2x_22 & IN2[48] | select_n2x_22 & (~ IN2[48]) | select_ne_22 & (~ IN2[49])  );
    wire logic pp_22_50;
    assign pp_22_50 = (select_e_22 & IN2[50] | select_2x_22 & IN2[49] | select_n2x_22 & (~ IN2[49]) | select_ne_22 & (~ IN2[50])  );
    wire logic pp_22_51;
    assign pp_22_51 = (select_e_22 & IN2[51] | select_2x_22 & IN2[50] | select_n2x_22 & (~ IN2[50]) | select_ne_22 & (~ IN2[51])  );
    wire logic pp_22_52;
    assign pp_22_52 = (select_e_22 & IN2[52] | select_2x_22 & IN2[51] | select_n2x_22 & (~ IN2[51]) | select_ne_22 & (~ IN2[52])  );
    wire logic pp_22_53;
    assign pp_22_53 = (select_e_22 & IN2[53] | select_2x_22 & IN2[52] | select_n2x_22 & (~ IN2[52]) | select_ne_22 & (~ IN2[53])  );
    wire logic pp_22_54;
    assign pp_22_54 = (select_e_22 & IN2[54] | select_2x_22 & IN2[53] | select_n2x_22 & (~ IN2[53]) | select_ne_22 & (~ IN2[54])  );
    wire logic pp_22_55;
    assign pp_22_55 = (select_e_22 & IN2[55] | select_2x_22 & IN2[54] | select_n2x_22 & (~ IN2[54]) | select_ne_22 & (~ IN2[55])  );
    wire logic pp_22_56;
    assign pp_22_56 = (select_e_22 & IN2[56] | select_2x_22 & IN2[55] | select_n2x_22 & (~ IN2[55]) | select_ne_22 & (~ IN2[56])  );
    wire logic pp_22_57;
    assign pp_22_57 = (select_e_22 & IN2[57] | select_2x_22 & IN2[56] | select_n2x_22 & (~ IN2[56]) | select_ne_22 & (~ IN2[57])  );
    wire logic pp_22_58;
    assign pp_22_58 = (select_e_22 & IN2[58] | select_2x_22 & IN2[57] | select_n2x_22 & (~ IN2[57]) | select_ne_22 & (~ IN2[58])  );
    wire logic pp_22_59;
    assign pp_22_59 = (select_e_22 & IN2[59] | select_2x_22 & IN2[58] | select_n2x_22 & (~ IN2[58]) | select_ne_22 & (~ IN2[59])  );
    wire logic pp_22_60;
    assign pp_22_60 = (select_e_22 & IN2[60] | select_2x_22 & IN2[59] | select_n2x_22 & (~ IN2[59]) | select_ne_22 & (~ IN2[60])  );
    wire logic pp_22_61;
    assign pp_22_61 = (select_e_22 & IN2[61] | select_2x_22 & IN2[60] | select_n2x_22 & (~ IN2[60]) | select_ne_22 & (~ IN2[61])  );
    wire logic pp_22_62;
    assign pp_22_62 = (select_e_22 & IN2[62] | select_2x_22 & IN2[61] | select_n2x_22 & (~ IN2[61]) | select_ne_22 & (~ IN2[62])  );
    wire logic pp_22_63;
    assign pp_22_63 = (select_e_22 & IN2[63] | select_2x_22 & IN2[62] | select_n2x_22 & (~ IN2[62]) | select_ne_22 & (~ IN2[63])  );
    wire logic pp_22_64;
    assign pp_22_64 = (select_e_22 & IN2[63] | select_2x_22 & IN2[63] | select_n2x_22 & (~ IN2[63]) | select_ne_22 & (~ IN2[63])  );
    wire logic pp_22_65;
    assign pp_22_65 = ~ (select_e_22 & IN2[63] | select_2x_22 & IN2[63] | select_n2x_22 & (~ IN2[63]) | select_ne_22 & (~ IN2[63])  );
    assign tcomp22 = select_ne_22 | select_n2x_22;
    
    // Signed Booth Radix-4 Partial Products Row 24
    wire logic select_e_23, select_ne_23, select_2x_23, tcomp23, select_n2x_23;
    assign select_e_23 = ((~ IN1[47]) & (IN1[46] ^ IN1[45]));
    assign select_ne_23 = IN1[47] &  (IN1[46] ^ IN1[45]);
    assign select_2x_23 = (~ IN1[47]) & IN1[46] & IN1[45];
    assign select_n2x_23 = IN1[47] & (~ IN1[46]) & (~ IN1[45]);
    wire logic pp_23_0;
    assign pp_23_0 = (select_e_23 & IN2[0] | select_2x_23 & 1'b0 | select_n2x_23 & 1'b1 | select_ne_23 & (~ IN2[0])  );
    wire logic pp_23_1;
    assign pp_23_1 = (select_e_23 & IN2[1] | select_2x_23 & IN2[0] | select_n2x_23 & (~ IN2[0]) | select_ne_23 & (~ IN2[1])  );
    wire logic pp_23_2;
    assign pp_23_2 = (select_e_23 & IN2[2] | select_2x_23 & IN2[1] | select_n2x_23 & (~ IN2[1]) | select_ne_23 & (~ IN2[2])  );
    wire logic pp_23_3;
    assign pp_23_3 = (select_e_23 & IN2[3] | select_2x_23 & IN2[2] | select_n2x_23 & (~ IN2[2]) | select_ne_23 & (~ IN2[3])  );
    wire logic pp_23_4;
    assign pp_23_4 = (select_e_23 & IN2[4] | select_2x_23 & IN2[3] | select_n2x_23 & (~ IN2[3]) | select_ne_23 & (~ IN2[4])  );
    wire logic pp_23_5;
    assign pp_23_5 = (select_e_23 & IN2[5] | select_2x_23 & IN2[4] | select_n2x_23 & (~ IN2[4]) | select_ne_23 & (~ IN2[5])  );
    wire logic pp_23_6;
    assign pp_23_6 = (select_e_23 & IN2[6] | select_2x_23 & IN2[5] | select_n2x_23 & (~ IN2[5]) | select_ne_23 & (~ IN2[6])  );
    wire logic pp_23_7;
    assign pp_23_7 = (select_e_23 & IN2[7] | select_2x_23 & IN2[6] | select_n2x_23 & (~ IN2[6]) | select_ne_23 & (~ IN2[7])  );
    wire logic pp_23_8;
    assign pp_23_8 = (select_e_23 & IN2[8] | select_2x_23 & IN2[7] | select_n2x_23 & (~ IN2[7]) | select_ne_23 & (~ IN2[8])  );
    wire logic pp_23_9;
    assign pp_23_9 = (select_e_23 & IN2[9] | select_2x_23 & IN2[8] | select_n2x_23 & (~ IN2[8]) | select_ne_23 & (~ IN2[9])  );
    wire logic pp_23_10;
    assign pp_23_10 = (select_e_23 & IN2[10] | select_2x_23 & IN2[9] | select_n2x_23 & (~ IN2[9]) | select_ne_23 & (~ IN2[10])  );
    wire logic pp_23_11;
    assign pp_23_11 = (select_e_23 & IN2[11] | select_2x_23 & IN2[10] | select_n2x_23 & (~ IN2[10]) | select_ne_23 & (~ IN2[11])  );
    wire logic pp_23_12;
    assign pp_23_12 = (select_e_23 & IN2[12] | select_2x_23 & IN2[11] | select_n2x_23 & (~ IN2[11]) | select_ne_23 & (~ IN2[12])  );
    wire logic pp_23_13;
    assign pp_23_13 = (select_e_23 & IN2[13] | select_2x_23 & IN2[12] | select_n2x_23 & (~ IN2[12]) | select_ne_23 & (~ IN2[13])  );
    wire logic pp_23_14;
    assign pp_23_14 = (select_e_23 & IN2[14] | select_2x_23 & IN2[13] | select_n2x_23 & (~ IN2[13]) | select_ne_23 & (~ IN2[14])  );
    wire logic pp_23_15;
    assign pp_23_15 = (select_e_23 & IN2[15] | select_2x_23 & IN2[14] | select_n2x_23 & (~ IN2[14]) | select_ne_23 & (~ IN2[15])  );
    wire logic pp_23_16;
    assign pp_23_16 = (select_e_23 & IN2[16] | select_2x_23 & IN2[15] | select_n2x_23 & (~ IN2[15]) | select_ne_23 & (~ IN2[16])  );
    wire logic pp_23_17;
    assign pp_23_17 = (select_e_23 & IN2[17] | select_2x_23 & IN2[16] | select_n2x_23 & (~ IN2[16]) | select_ne_23 & (~ IN2[17])  );
    wire logic pp_23_18;
    assign pp_23_18 = (select_e_23 & IN2[18] | select_2x_23 & IN2[17] | select_n2x_23 & (~ IN2[17]) | select_ne_23 & (~ IN2[18])  );
    wire logic pp_23_19;
    assign pp_23_19 = (select_e_23 & IN2[19] | select_2x_23 & IN2[18] | select_n2x_23 & (~ IN2[18]) | select_ne_23 & (~ IN2[19])  );
    wire logic pp_23_20;
    assign pp_23_20 = (select_e_23 & IN2[20] | select_2x_23 & IN2[19] | select_n2x_23 & (~ IN2[19]) | select_ne_23 & (~ IN2[20])  );
    wire logic pp_23_21;
    assign pp_23_21 = (select_e_23 & IN2[21] | select_2x_23 & IN2[20] | select_n2x_23 & (~ IN2[20]) | select_ne_23 & (~ IN2[21])  );
    wire logic pp_23_22;
    assign pp_23_22 = (select_e_23 & IN2[22] | select_2x_23 & IN2[21] | select_n2x_23 & (~ IN2[21]) | select_ne_23 & (~ IN2[22])  );
    wire logic pp_23_23;
    assign pp_23_23 = (select_e_23 & IN2[23] | select_2x_23 & IN2[22] | select_n2x_23 & (~ IN2[22]) | select_ne_23 & (~ IN2[23])  );
    wire logic pp_23_24;
    assign pp_23_24 = (select_e_23 & IN2[24] | select_2x_23 & IN2[23] | select_n2x_23 & (~ IN2[23]) | select_ne_23 & (~ IN2[24])  );
    wire logic pp_23_25;
    assign pp_23_25 = (select_e_23 & IN2[25] | select_2x_23 & IN2[24] | select_n2x_23 & (~ IN2[24]) | select_ne_23 & (~ IN2[25])  );
    wire logic pp_23_26;
    assign pp_23_26 = (select_e_23 & IN2[26] | select_2x_23 & IN2[25] | select_n2x_23 & (~ IN2[25]) | select_ne_23 & (~ IN2[26])  );
    wire logic pp_23_27;
    assign pp_23_27 = (select_e_23 & IN2[27] | select_2x_23 & IN2[26] | select_n2x_23 & (~ IN2[26]) | select_ne_23 & (~ IN2[27])  );
    wire logic pp_23_28;
    assign pp_23_28 = (select_e_23 & IN2[28] | select_2x_23 & IN2[27] | select_n2x_23 & (~ IN2[27]) | select_ne_23 & (~ IN2[28])  );
    wire logic pp_23_29;
    assign pp_23_29 = (select_e_23 & IN2[29] | select_2x_23 & IN2[28] | select_n2x_23 & (~ IN2[28]) | select_ne_23 & (~ IN2[29])  );
    wire logic pp_23_30;
    assign pp_23_30 = (select_e_23 & IN2[30] | select_2x_23 & IN2[29] | select_n2x_23 & (~ IN2[29]) | select_ne_23 & (~ IN2[30])  );
    wire logic pp_23_31;
    assign pp_23_31 = (select_e_23 & IN2[31] | select_2x_23 & IN2[30] | select_n2x_23 & (~ IN2[30]) | select_ne_23 & (~ IN2[31])  );
    wire logic pp_23_32;
    assign pp_23_32 = (select_e_23 & IN2[32] | select_2x_23 & IN2[31] | select_n2x_23 & (~ IN2[31]) | select_ne_23 & (~ IN2[32])  );
    wire logic pp_23_33;
    assign pp_23_33 = (select_e_23 & IN2[33] | select_2x_23 & IN2[32] | select_n2x_23 & (~ IN2[32]) | select_ne_23 & (~ IN2[33])  );
    wire logic pp_23_34;
    assign pp_23_34 = (select_e_23 & IN2[34] | select_2x_23 & IN2[33] | select_n2x_23 & (~ IN2[33]) | select_ne_23 & (~ IN2[34])  );
    wire logic pp_23_35;
    assign pp_23_35 = (select_e_23 & IN2[35] | select_2x_23 & IN2[34] | select_n2x_23 & (~ IN2[34]) | select_ne_23 & (~ IN2[35])  );
    wire logic pp_23_36;
    assign pp_23_36 = (select_e_23 & IN2[36] | select_2x_23 & IN2[35] | select_n2x_23 & (~ IN2[35]) | select_ne_23 & (~ IN2[36])  );
    wire logic pp_23_37;
    assign pp_23_37 = (select_e_23 & IN2[37] | select_2x_23 & IN2[36] | select_n2x_23 & (~ IN2[36]) | select_ne_23 & (~ IN2[37])  );
    wire logic pp_23_38;
    assign pp_23_38 = (select_e_23 & IN2[38] | select_2x_23 & IN2[37] | select_n2x_23 & (~ IN2[37]) | select_ne_23 & (~ IN2[38])  );
    wire logic pp_23_39;
    assign pp_23_39 = (select_e_23 & IN2[39] | select_2x_23 & IN2[38] | select_n2x_23 & (~ IN2[38]) | select_ne_23 & (~ IN2[39])  );
    wire logic pp_23_40;
    assign pp_23_40 = (select_e_23 & IN2[40] | select_2x_23 & IN2[39] | select_n2x_23 & (~ IN2[39]) | select_ne_23 & (~ IN2[40])  );
    wire logic pp_23_41;
    assign pp_23_41 = (select_e_23 & IN2[41] | select_2x_23 & IN2[40] | select_n2x_23 & (~ IN2[40]) | select_ne_23 & (~ IN2[41])  );
    wire logic pp_23_42;
    assign pp_23_42 = (select_e_23 & IN2[42] | select_2x_23 & IN2[41] | select_n2x_23 & (~ IN2[41]) | select_ne_23 & (~ IN2[42])  );
    wire logic pp_23_43;
    assign pp_23_43 = (select_e_23 & IN2[43] | select_2x_23 & IN2[42] | select_n2x_23 & (~ IN2[42]) | select_ne_23 & (~ IN2[43])  );
    wire logic pp_23_44;
    assign pp_23_44 = (select_e_23 & IN2[44] | select_2x_23 & IN2[43] | select_n2x_23 & (~ IN2[43]) | select_ne_23 & (~ IN2[44])  );
    wire logic pp_23_45;
    assign pp_23_45 = (select_e_23 & IN2[45] | select_2x_23 & IN2[44] | select_n2x_23 & (~ IN2[44]) | select_ne_23 & (~ IN2[45])  );
    wire logic pp_23_46;
    assign pp_23_46 = (select_e_23 & IN2[46] | select_2x_23 & IN2[45] | select_n2x_23 & (~ IN2[45]) | select_ne_23 & (~ IN2[46])  );
    wire logic pp_23_47;
    assign pp_23_47 = (select_e_23 & IN2[47] | select_2x_23 & IN2[46] | select_n2x_23 & (~ IN2[46]) | select_ne_23 & (~ IN2[47])  );
    wire logic pp_23_48;
    assign pp_23_48 = (select_e_23 & IN2[48] | select_2x_23 & IN2[47] | select_n2x_23 & (~ IN2[47]) | select_ne_23 & (~ IN2[48])  );
    wire logic pp_23_49;
    assign pp_23_49 = (select_e_23 & IN2[49] | select_2x_23 & IN2[48] | select_n2x_23 & (~ IN2[48]) | select_ne_23 & (~ IN2[49])  );
    wire logic pp_23_50;
    assign pp_23_50 = (select_e_23 & IN2[50] | select_2x_23 & IN2[49] | select_n2x_23 & (~ IN2[49]) | select_ne_23 & (~ IN2[50])  );
    wire logic pp_23_51;
    assign pp_23_51 = (select_e_23 & IN2[51] | select_2x_23 & IN2[50] | select_n2x_23 & (~ IN2[50]) | select_ne_23 & (~ IN2[51])  );
    wire logic pp_23_52;
    assign pp_23_52 = (select_e_23 & IN2[52] | select_2x_23 & IN2[51] | select_n2x_23 & (~ IN2[51]) | select_ne_23 & (~ IN2[52])  );
    wire logic pp_23_53;
    assign pp_23_53 = (select_e_23 & IN2[53] | select_2x_23 & IN2[52] | select_n2x_23 & (~ IN2[52]) | select_ne_23 & (~ IN2[53])  );
    wire logic pp_23_54;
    assign pp_23_54 = (select_e_23 & IN2[54] | select_2x_23 & IN2[53] | select_n2x_23 & (~ IN2[53]) | select_ne_23 & (~ IN2[54])  );
    wire logic pp_23_55;
    assign pp_23_55 = (select_e_23 & IN2[55] | select_2x_23 & IN2[54] | select_n2x_23 & (~ IN2[54]) | select_ne_23 & (~ IN2[55])  );
    wire logic pp_23_56;
    assign pp_23_56 = (select_e_23 & IN2[56] | select_2x_23 & IN2[55] | select_n2x_23 & (~ IN2[55]) | select_ne_23 & (~ IN2[56])  );
    wire logic pp_23_57;
    assign pp_23_57 = (select_e_23 & IN2[57] | select_2x_23 & IN2[56] | select_n2x_23 & (~ IN2[56]) | select_ne_23 & (~ IN2[57])  );
    wire logic pp_23_58;
    assign pp_23_58 = (select_e_23 & IN2[58] | select_2x_23 & IN2[57] | select_n2x_23 & (~ IN2[57]) | select_ne_23 & (~ IN2[58])  );
    wire logic pp_23_59;
    assign pp_23_59 = (select_e_23 & IN2[59] | select_2x_23 & IN2[58] | select_n2x_23 & (~ IN2[58]) | select_ne_23 & (~ IN2[59])  );
    wire logic pp_23_60;
    assign pp_23_60 = (select_e_23 & IN2[60] | select_2x_23 & IN2[59] | select_n2x_23 & (~ IN2[59]) | select_ne_23 & (~ IN2[60])  );
    wire logic pp_23_61;
    assign pp_23_61 = (select_e_23 & IN2[61] | select_2x_23 & IN2[60] | select_n2x_23 & (~ IN2[60]) | select_ne_23 & (~ IN2[61])  );
    wire logic pp_23_62;
    assign pp_23_62 = (select_e_23 & IN2[62] | select_2x_23 & IN2[61] | select_n2x_23 & (~ IN2[61]) | select_ne_23 & (~ IN2[62])  );
    wire logic pp_23_63;
    assign pp_23_63 = (select_e_23 & IN2[63] | select_2x_23 & IN2[62] | select_n2x_23 & (~ IN2[62]) | select_ne_23 & (~ IN2[63])  );
    wire logic pp_23_64;
    assign pp_23_64 = (select_e_23 & IN2[63] | select_2x_23 & IN2[63] | select_n2x_23 & (~ IN2[63]) | select_ne_23 & (~ IN2[63])  );
    wire logic pp_23_65;
    assign pp_23_65 = ~ (select_e_23 & IN2[63] | select_2x_23 & IN2[63] | select_n2x_23 & (~ IN2[63]) | select_ne_23 & (~ IN2[63])  );
    assign tcomp23 = select_ne_23 | select_n2x_23;
    
    // Signed Booth Radix-4 Partial Products Row 25
    wire logic select_e_24, select_ne_24, select_2x_24, tcomp24, select_n2x_24;
    assign select_e_24 = ((~ IN1[49]) & (IN1[48] ^ IN1[47]));
    assign select_ne_24 = IN1[49] &  (IN1[48] ^ IN1[47]);
    assign select_2x_24 = (~ IN1[49]) & IN1[48] & IN1[47];
    assign select_n2x_24 = IN1[49] & (~ IN1[48]) & (~ IN1[47]);
    wire logic pp_24_0;
    assign pp_24_0 = (select_e_24 & IN2[0] | select_2x_24 & 1'b0 | select_n2x_24 & 1'b1 | select_ne_24 & (~ IN2[0])  );
    wire logic pp_24_1;
    assign pp_24_1 = (select_e_24 & IN2[1] | select_2x_24 & IN2[0] | select_n2x_24 & (~ IN2[0]) | select_ne_24 & (~ IN2[1])  );
    wire logic pp_24_2;
    assign pp_24_2 = (select_e_24 & IN2[2] | select_2x_24 & IN2[1] | select_n2x_24 & (~ IN2[1]) | select_ne_24 & (~ IN2[2])  );
    wire logic pp_24_3;
    assign pp_24_3 = (select_e_24 & IN2[3] | select_2x_24 & IN2[2] | select_n2x_24 & (~ IN2[2]) | select_ne_24 & (~ IN2[3])  );
    wire logic pp_24_4;
    assign pp_24_4 = (select_e_24 & IN2[4] | select_2x_24 & IN2[3] | select_n2x_24 & (~ IN2[3]) | select_ne_24 & (~ IN2[4])  );
    wire logic pp_24_5;
    assign pp_24_5 = (select_e_24 & IN2[5] | select_2x_24 & IN2[4] | select_n2x_24 & (~ IN2[4]) | select_ne_24 & (~ IN2[5])  );
    wire logic pp_24_6;
    assign pp_24_6 = (select_e_24 & IN2[6] | select_2x_24 & IN2[5] | select_n2x_24 & (~ IN2[5]) | select_ne_24 & (~ IN2[6])  );
    wire logic pp_24_7;
    assign pp_24_7 = (select_e_24 & IN2[7] | select_2x_24 & IN2[6] | select_n2x_24 & (~ IN2[6]) | select_ne_24 & (~ IN2[7])  );
    wire logic pp_24_8;
    assign pp_24_8 = (select_e_24 & IN2[8] | select_2x_24 & IN2[7] | select_n2x_24 & (~ IN2[7]) | select_ne_24 & (~ IN2[8])  );
    wire logic pp_24_9;
    assign pp_24_9 = (select_e_24 & IN2[9] | select_2x_24 & IN2[8] | select_n2x_24 & (~ IN2[8]) | select_ne_24 & (~ IN2[9])  );
    wire logic pp_24_10;
    assign pp_24_10 = (select_e_24 & IN2[10] | select_2x_24 & IN2[9] | select_n2x_24 & (~ IN2[9]) | select_ne_24 & (~ IN2[10])  );
    wire logic pp_24_11;
    assign pp_24_11 = (select_e_24 & IN2[11] | select_2x_24 & IN2[10] | select_n2x_24 & (~ IN2[10]) | select_ne_24 & (~ IN2[11])  );
    wire logic pp_24_12;
    assign pp_24_12 = (select_e_24 & IN2[12] | select_2x_24 & IN2[11] | select_n2x_24 & (~ IN2[11]) | select_ne_24 & (~ IN2[12])  );
    wire logic pp_24_13;
    assign pp_24_13 = (select_e_24 & IN2[13] | select_2x_24 & IN2[12] | select_n2x_24 & (~ IN2[12]) | select_ne_24 & (~ IN2[13])  );
    wire logic pp_24_14;
    assign pp_24_14 = (select_e_24 & IN2[14] | select_2x_24 & IN2[13] | select_n2x_24 & (~ IN2[13]) | select_ne_24 & (~ IN2[14])  );
    wire logic pp_24_15;
    assign pp_24_15 = (select_e_24 & IN2[15] | select_2x_24 & IN2[14] | select_n2x_24 & (~ IN2[14]) | select_ne_24 & (~ IN2[15])  );
    wire logic pp_24_16;
    assign pp_24_16 = (select_e_24 & IN2[16] | select_2x_24 & IN2[15] | select_n2x_24 & (~ IN2[15]) | select_ne_24 & (~ IN2[16])  );
    wire logic pp_24_17;
    assign pp_24_17 = (select_e_24 & IN2[17] | select_2x_24 & IN2[16] | select_n2x_24 & (~ IN2[16]) | select_ne_24 & (~ IN2[17])  );
    wire logic pp_24_18;
    assign pp_24_18 = (select_e_24 & IN2[18] | select_2x_24 & IN2[17] | select_n2x_24 & (~ IN2[17]) | select_ne_24 & (~ IN2[18])  );
    wire logic pp_24_19;
    assign pp_24_19 = (select_e_24 & IN2[19] | select_2x_24 & IN2[18] | select_n2x_24 & (~ IN2[18]) | select_ne_24 & (~ IN2[19])  );
    wire logic pp_24_20;
    assign pp_24_20 = (select_e_24 & IN2[20] | select_2x_24 & IN2[19] | select_n2x_24 & (~ IN2[19]) | select_ne_24 & (~ IN2[20])  );
    wire logic pp_24_21;
    assign pp_24_21 = (select_e_24 & IN2[21] | select_2x_24 & IN2[20] | select_n2x_24 & (~ IN2[20]) | select_ne_24 & (~ IN2[21])  );
    wire logic pp_24_22;
    assign pp_24_22 = (select_e_24 & IN2[22] | select_2x_24 & IN2[21] | select_n2x_24 & (~ IN2[21]) | select_ne_24 & (~ IN2[22])  );
    wire logic pp_24_23;
    assign pp_24_23 = (select_e_24 & IN2[23] | select_2x_24 & IN2[22] | select_n2x_24 & (~ IN2[22]) | select_ne_24 & (~ IN2[23])  );
    wire logic pp_24_24;
    assign pp_24_24 = (select_e_24 & IN2[24] | select_2x_24 & IN2[23] | select_n2x_24 & (~ IN2[23]) | select_ne_24 & (~ IN2[24])  );
    wire logic pp_24_25;
    assign pp_24_25 = (select_e_24 & IN2[25] | select_2x_24 & IN2[24] | select_n2x_24 & (~ IN2[24]) | select_ne_24 & (~ IN2[25])  );
    wire logic pp_24_26;
    assign pp_24_26 = (select_e_24 & IN2[26] | select_2x_24 & IN2[25] | select_n2x_24 & (~ IN2[25]) | select_ne_24 & (~ IN2[26])  );
    wire logic pp_24_27;
    assign pp_24_27 = (select_e_24 & IN2[27] | select_2x_24 & IN2[26] | select_n2x_24 & (~ IN2[26]) | select_ne_24 & (~ IN2[27])  );
    wire logic pp_24_28;
    assign pp_24_28 = (select_e_24 & IN2[28] | select_2x_24 & IN2[27] | select_n2x_24 & (~ IN2[27]) | select_ne_24 & (~ IN2[28])  );
    wire logic pp_24_29;
    assign pp_24_29 = (select_e_24 & IN2[29] | select_2x_24 & IN2[28] | select_n2x_24 & (~ IN2[28]) | select_ne_24 & (~ IN2[29])  );
    wire logic pp_24_30;
    assign pp_24_30 = (select_e_24 & IN2[30] | select_2x_24 & IN2[29] | select_n2x_24 & (~ IN2[29]) | select_ne_24 & (~ IN2[30])  );
    wire logic pp_24_31;
    assign pp_24_31 = (select_e_24 & IN2[31] | select_2x_24 & IN2[30] | select_n2x_24 & (~ IN2[30]) | select_ne_24 & (~ IN2[31])  );
    wire logic pp_24_32;
    assign pp_24_32 = (select_e_24 & IN2[32] | select_2x_24 & IN2[31] | select_n2x_24 & (~ IN2[31]) | select_ne_24 & (~ IN2[32])  );
    wire logic pp_24_33;
    assign pp_24_33 = (select_e_24 & IN2[33] | select_2x_24 & IN2[32] | select_n2x_24 & (~ IN2[32]) | select_ne_24 & (~ IN2[33])  );
    wire logic pp_24_34;
    assign pp_24_34 = (select_e_24 & IN2[34] | select_2x_24 & IN2[33] | select_n2x_24 & (~ IN2[33]) | select_ne_24 & (~ IN2[34])  );
    wire logic pp_24_35;
    assign pp_24_35 = (select_e_24 & IN2[35] | select_2x_24 & IN2[34] | select_n2x_24 & (~ IN2[34]) | select_ne_24 & (~ IN2[35])  );
    wire logic pp_24_36;
    assign pp_24_36 = (select_e_24 & IN2[36] | select_2x_24 & IN2[35] | select_n2x_24 & (~ IN2[35]) | select_ne_24 & (~ IN2[36])  );
    wire logic pp_24_37;
    assign pp_24_37 = (select_e_24 & IN2[37] | select_2x_24 & IN2[36] | select_n2x_24 & (~ IN2[36]) | select_ne_24 & (~ IN2[37])  );
    wire logic pp_24_38;
    assign pp_24_38 = (select_e_24 & IN2[38] | select_2x_24 & IN2[37] | select_n2x_24 & (~ IN2[37]) | select_ne_24 & (~ IN2[38])  );
    wire logic pp_24_39;
    assign pp_24_39 = (select_e_24 & IN2[39] | select_2x_24 & IN2[38] | select_n2x_24 & (~ IN2[38]) | select_ne_24 & (~ IN2[39])  );
    wire logic pp_24_40;
    assign pp_24_40 = (select_e_24 & IN2[40] | select_2x_24 & IN2[39] | select_n2x_24 & (~ IN2[39]) | select_ne_24 & (~ IN2[40])  );
    wire logic pp_24_41;
    assign pp_24_41 = (select_e_24 & IN2[41] | select_2x_24 & IN2[40] | select_n2x_24 & (~ IN2[40]) | select_ne_24 & (~ IN2[41])  );
    wire logic pp_24_42;
    assign pp_24_42 = (select_e_24 & IN2[42] | select_2x_24 & IN2[41] | select_n2x_24 & (~ IN2[41]) | select_ne_24 & (~ IN2[42])  );
    wire logic pp_24_43;
    assign pp_24_43 = (select_e_24 & IN2[43] | select_2x_24 & IN2[42] | select_n2x_24 & (~ IN2[42]) | select_ne_24 & (~ IN2[43])  );
    wire logic pp_24_44;
    assign pp_24_44 = (select_e_24 & IN2[44] | select_2x_24 & IN2[43] | select_n2x_24 & (~ IN2[43]) | select_ne_24 & (~ IN2[44])  );
    wire logic pp_24_45;
    assign pp_24_45 = (select_e_24 & IN2[45] | select_2x_24 & IN2[44] | select_n2x_24 & (~ IN2[44]) | select_ne_24 & (~ IN2[45])  );
    wire logic pp_24_46;
    assign pp_24_46 = (select_e_24 & IN2[46] | select_2x_24 & IN2[45] | select_n2x_24 & (~ IN2[45]) | select_ne_24 & (~ IN2[46])  );
    wire logic pp_24_47;
    assign pp_24_47 = (select_e_24 & IN2[47] | select_2x_24 & IN2[46] | select_n2x_24 & (~ IN2[46]) | select_ne_24 & (~ IN2[47])  );
    wire logic pp_24_48;
    assign pp_24_48 = (select_e_24 & IN2[48] | select_2x_24 & IN2[47] | select_n2x_24 & (~ IN2[47]) | select_ne_24 & (~ IN2[48])  );
    wire logic pp_24_49;
    assign pp_24_49 = (select_e_24 & IN2[49] | select_2x_24 & IN2[48] | select_n2x_24 & (~ IN2[48]) | select_ne_24 & (~ IN2[49])  );
    wire logic pp_24_50;
    assign pp_24_50 = (select_e_24 & IN2[50] | select_2x_24 & IN2[49] | select_n2x_24 & (~ IN2[49]) | select_ne_24 & (~ IN2[50])  );
    wire logic pp_24_51;
    assign pp_24_51 = (select_e_24 & IN2[51] | select_2x_24 & IN2[50] | select_n2x_24 & (~ IN2[50]) | select_ne_24 & (~ IN2[51])  );
    wire logic pp_24_52;
    assign pp_24_52 = (select_e_24 & IN2[52] | select_2x_24 & IN2[51] | select_n2x_24 & (~ IN2[51]) | select_ne_24 & (~ IN2[52])  );
    wire logic pp_24_53;
    assign pp_24_53 = (select_e_24 & IN2[53] | select_2x_24 & IN2[52] | select_n2x_24 & (~ IN2[52]) | select_ne_24 & (~ IN2[53])  );
    wire logic pp_24_54;
    assign pp_24_54 = (select_e_24 & IN2[54] | select_2x_24 & IN2[53] | select_n2x_24 & (~ IN2[53]) | select_ne_24 & (~ IN2[54])  );
    wire logic pp_24_55;
    assign pp_24_55 = (select_e_24 & IN2[55] | select_2x_24 & IN2[54] | select_n2x_24 & (~ IN2[54]) | select_ne_24 & (~ IN2[55])  );
    wire logic pp_24_56;
    assign pp_24_56 = (select_e_24 & IN2[56] | select_2x_24 & IN2[55] | select_n2x_24 & (~ IN2[55]) | select_ne_24 & (~ IN2[56])  );
    wire logic pp_24_57;
    assign pp_24_57 = (select_e_24 & IN2[57] | select_2x_24 & IN2[56] | select_n2x_24 & (~ IN2[56]) | select_ne_24 & (~ IN2[57])  );
    wire logic pp_24_58;
    assign pp_24_58 = (select_e_24 & IN2[58] | select_2x_24 & IN2[57] | select_n2x_24 & (~ IN2[57]) | select_ne_24 & (~ IN2[58])  );
    wire logic pp_24_59;
    assign pp_24_59 = (select_e_24 & IN2[59] | select_2x_24 & IN2[58] | select_n2x_24 & (~ IN2[58]) | select_ne_24 & (~ IN2[59])  );
    wire logic pp_24_60;
    assign pp_24_60 = (select_e_24 & IN2[60] | select_2x_24 & IN2[59] | select_n2x_24 & (~ IN2[59]) | select_ne_24 & (~ IN2[60])  );
    wire logic pp_24_61;
    assign pp_24_61 = (select_e_24 & IN2[61] | select_2x_24 & IN2[60] | select_n2x_24 & (~ IN2[60]) | select_ne_24 & (~ IN2[61])  );
    wire logic pp_24_62;
    assign pp_24_62 = (select_e_24 & IN2[62] | select_2x_24 & IN2[61] | select_n2x_24 & (~ IN2[61]) | select_ne_24 & (~ IN2[62])  );
    wire logic pp_24_63;
    assign pp_24_63 = (select_e_24 & IN2[63] | select_2x_24 & IN2[62] | select_n2x_24 & (~ IN2[62]) | select_ne_24 & (~ IN2[63])  );
    wire logic pp_24_64;
    assign pp_24_64 = (select_e_24 & IN2[63] | select_2x_24 & IN2[63] | select_n2x_24 & (~ IN2[63]) | select_ne_24 & (~ IN2[63])  );
    wire logic pp_24_65;
    assign pp_24_65 = ~ (select_e_24 & IN2[63] | select_2x_24 & IN2[63] | select_n2x_24 & (~ IN2[63]) | select_ne_24 & (~ IN2[63])  );
    assign tcomp24 = select_ne_24 | select_n2x_24;
    
    // Signed Booth Radix-4 Partial Products Row 26
    wire logic select_e_25, select_ne_25, select_2x_25, tcomp25, select_n2x_25;
    assign select_e_25 = ((~ IN1[51]) & (IN1[50] ^ IN1[49]));
    assign select_ne_25 = IN1[51] &  (IN1[50] ^ IN1[49]);
    assign select_2x_25 = (~ IN1[51]) & IN1[50] & IN1[49];
    assign select_n2x_25 = IN1[51] & (~ IN1[50]) & (~ IN1[49]);
    wire logic pp_25_0;
    assign pp_25_0 = (select_e_25 & IN2[0] | select_2x_25 & 1'b0 | select_n2x_25 & 1'b1 | select_ne_25 & (~ IN2[0])  );
    wire logic pp_25_1;
    assign pp_25_1 = (select_e_25 & IN2[1] | select_2x_25 & IN2[0] | select_n2x_25 & (~ IN2[0]) | select_ne_25 & (~ IN2[1])  );
    wire logic pp_25_2;
    assign pp_25_2 = (select_e_25 & IN2[2] | select_2x_25 & IN2[1] | select_n2x_25 & (~ IN2[1]) | select_ne_25 & (~ IN2[2])  );
    wire logic pp_25_3;
    assign pp_25_3 = (select_e_25 & IN2[3] | select_2x_25 & IN2[2] | select_n2x_25 & (~ IN2[2]) | select_ne_25 & (~ IN2[3])  );
    wire logic pp_25_4;
    assign pp_25_4 = (select_e_25 & IN2[4] | select_2x_25 & IN2[3] | select_n2x_25 & (~ IN2[3]) | select_ne_25 & (~ IN2[4])  );
    wire logic pp_25_5;
    assign pp_25_5 = (select_e_25 & IN2[5] | select_2x_25 & IN2[4] | select_n2x_25 & (~ IN2[4]) | select_ne_25 & (~ IN2[5])  );
    wire logic pp_25_6;
    assign pp_25_6 = (select_e_25 & IN2[6] | select_2x_25 & IN2[5] | select_n2x_25 & (~ IN2[5]) | select_ne_25 & (~ IN2[6])  );
    wire logic pp_25_7;
    assign pp_25_7 = (select_e_25 & IN2[7] | select_2x_25 & IN2[6] | select_n2x_25 & (~ IN2[6]) | select_ne_25 & (~ IN2[7])  );
    wire logic pp_25_8;
    assign pp_25_8 = (select_e_25 & IN2[8] | select_2x_25 & IN2[7] | select_n2x_25 & (~ IN2[7]) | select_ne_25 & (~ IN2[8])  );
    wire logic pp_25_9;
    assign pp_25_9 = (select_e_25 & IN2[9] | select_2x_25 & IN2[8] | select_n2x_25 & (~ IN2[8]) | select_ne_25 & (~ IN2[9])  );
    wire logic pp_25_10;
    assign pp_25_10 = (select_e_25 & IN2[10] | select_2x_25 & IN2[9] | select_n2x_25 & (~ IN2[9]) | select_ne_25 & (~ IN2[10])  );
    wire logic pp_25_11;
    assign pp_25_11 = (select_e_25 & IN2[11] | select_2x_25 & IN2[10] | select_n2x_25 & (~ IN2[10]) | select_ne_25 & (~ IN2[11])  );
    wire logic pp_25_12;
    assign pp_25_12 = (select_e_25 & IN2[12] | select_2x_25 & IN2[11] | select_n2x_25 & (~ IN2[11]) | select_ne_25 & (~ IN2[12])  );
    wire logic pp_25_13;
    assign pp_25_13 = (select_e_25 & IN2[13] | select_2x_25 & IN2[12] | select_n2x_25 & (~ IN2[12]) | select_ne_25 & (~ IN2[13])  );
    wire logic pp_25_14;
    assign pp_25_14 = (select_e_25 & IN2[14] | select_2x_25 & IN2[13] | select_n2x_25 & (~ IN2[13]) | select_ne_25 & (~ IN2[14])  );
    wire logic pp_25_15;
    assign pp_25_15 = (select_e_25 & IN2[15] | select_2x_25 & IN2[14] | select_n2x_25 & (~ IN2[14]) | select_ne_25 & (~ IN2[15])  );
    wire logic pp_25_16;
    assign pp_25_16 = (select_e_25 & IN2[16] | select_2x_25 & IN2[15] | select_n2x_25 & (~ IN2[15]) | select_ne_25 & (~ IN2[16])  );
    wire logic pp_25_17;
    assign pp_25_17 = (select_e_25 & IN2[17] | select_2x_25 & IN2[16] | select_n2x_25 & (~ IN2[16]) | select_ne_25 & (~ IN2[17])  );
    wire logic pp_25_18;
    assign pp_25_18 = (select_e_25 & IN2[18] | select_2x_25 & IN2[17] | select_n2x_25 & (~ IN2[17]) | select_ne_25 & (~ IN2[18])  );
    wire logic pp_25_19;
    assign pp_25_19 = (select_e_25 & IN2[19] | select_2x_25 & IN2[18] | select_n2x_25 & (~ IN2[18]) | select_ne_25 & (~ IN2[19])  );
    wire logic pp_25_20;
    assign pp_25_20 = (select_e_25 & IN2[20] | select_2x_25 & IN2[19] | select_n2x_25 & (~ IN2[19]) | select_ne_25 & (~ IN2[20])  );
    wire logic pp_25_21;
    assign pp_25_21 = (select_e_25 & IN2[21] | select_2x_25 & IN2[20] | select_n2x_25 & (~ IN2[20]) | select_ne_25 & (~ IN2[21])  );
    wire logic pp_25_22;
    assign pp_25_22 = (select_e_25 & IN2[22] | select_2x_25 & IN2[21] | select_n2x_25 & (~ IN2[21]) | select_ne_25 & (~ IN2[22])  );
    wire logic pp_25_23;
    assign pp_25_23 = (select_e_25 & IN2[23] | select_2x_25 & IN2[22] | select_n2x_25 & (~ IN2[22]) | select_ne_25 & (~ IN2[23])  );
    wire logic pp_25_24;
    assign pp_25_24 = (select_e_25 & IN2[24] | select_2x_25 & IN2[23] | select_n2x_25 & (~ IN2[23]) | select_ne_25 & (~ IN2[24])  );
    wire logic pp_25_25;
    assign pp_25_25 = (select_e_25 & IN2[25] | select_2x_25 & IN2[24] | select_n2x_25 & (~ IN2[24]) | select_ne_25 & (~ IN2[25])  );
    wire logic pp_25_26;
    assign pp_25_26 = (select_e_25 & IN2[26] | select_2x_25 & IN2[25] | select_n2x_25 & (~ IN2[25]) | select_ne_25 & (~ IN2[26])  );
    wire logic pp_25_27;
    assign pp_25_27 = (select_e_25 & IN2[27] | select_2x_25 & IN2[26] | select_n2x_25 & (~ IN2[26]) | select_ne_25 & (~ IN2[27])  );
    wire logic pp_25_28;
    assign pp_25_28 = (select_e_25 & IN2[28] | select_2x_25 & IN2[27] | select_n2x_25 & (~ IN2[27]) | select_ne_25 & (~ IN2[28])  );
    wire logic pp_25_29;
    assign pp_25_29 = (select_e_25 & IN2[29] | select_2x_25 & IN2[28] | select_n2x_25 & (~ IN2[28]) | select_ne_25 & (~ IN2[29])  );
    wire logic pp_25_30;
    assign pp_25_30 = (select_e_25 & IN2[30] | select_2x_25 & IN2[29] | select_n2x_25 & (~ IN2[29]) | select_ne_25 & (~ IN2[30])  );
    wire logic pp_25_31;
    assign pp_25_31 = (select_e_25 & IN2[31] | select_2x_25 & IN2[30] | select_n2x_25 & (~ IN2[30]) | select_ne_25 & (~ IN2[31])  );
    wire logic pp_25_32;
    assign pp_25_32 = (select_e_25 & IN2[32] | select_2x_25 & IN2[31] | select_n2x_25 & (~ IN2[31]) | select_ne_25 & (~ IN2[32])  );
    wire logic pp_25_33;
    assign pp_25_33 = (select_e_25 & IN2[33] | select_2x_25 & IN2[32] | select_n2x_25 & (~ IN2[32]) | select_ne_25 & (~ IN2[33])  );
    wire logic pp_25_34;
    assign pp_25_34 = (select_e_25 & IN2[34] | select_2x_25 & IN2[33] | select_n2x_25 & (~ IN2[33]) | select_ne_25 & (~ IN2[34])  );
    wire logic pp_25_35;
    assign pp_25_35 = (select_e_25 & IN2[35] | select_2x_25 & IN2[34] | select_n2x_25 & (~ IN2[34]) | select_ne_25 & (~ IN2[35])  );
    wire logic pp_25_36;
    assign pp_25_36 = (select_e_25 & IN2[36] | select_2x_25 & IN2[35] | select_n2x_25 & (~ IN2[35]) | select_ne_25 & (~ IN2[36])  );
    wire logic pp_25_37;
    assign pp_25_37 = (select_e_25 & IN2[37] | select_2x_25 & IN2[36] | select_n2x_25 & (~ IN2[36]) | select_ne_25 & (~ IN2[37])  );
    wire logic pp_25_38;
    assign pp_25_38 = (select_e_25 & IN2[38] | select_2x_25 & IN2[37] | select_n2x_25 & (~ IN2[37]) | select_ne_25 & (~ IN2[38])  );
    wire logic pp_25_39;
    assign pp_25_39 = (select_e_25 & IN2[39] | select_2x_25 & IN2[38] | select_n2x_25 & (~ IN2[38]) | select_ne_25 & (~ IN2[39])  );
    wire logic pp_25_40;
    assign pp_25_40 = (select_e_25 & IN2[40] | select_2x_25 & IN2[39] | select_n2x_25 & (~ IN2[39]) | select_ne_25 & (~ IN2[40])  );
    wire logic pp_25_41;
    assign pp_25_41 = (select_e_25 & IN2[41] | select_2x_25 & IN2[40] | select_n2x_25 & (~ IN2[40]) | select_ne_25 & (~ IN2[41])  );
    wire logic pp_25_42;
    assign pp_25_42 = (select_e_25 & IN2[42] | select_2x_25 & IN2[41] | select_n2x_25 & (~ IN2[41]) | select_ne_25 & (~ IN2[42])  );
    wire logic pp_25_43;
    assign pp_25_43 = (select_e_25 & IN2[43] | select_2x_25 & IN2[42] | select_n2x_25 & (~ IN2[42]) | select_ne_25 & (~ IN2[43])  );
    wire logic pp_25_44;
    assign pp_25_44 = (select_e_25 & IN2[44] | select_2x_25 & IN2[43] | select_n2x_25 & (~ IN2[43]) | select_ne_25 & (~ IN2[44])  );
    wire logic pp_25_45;
    assign pp_25_45 = (select_e_25 & IN2[45] | select_2x_25 & IN2[44] | select_n2x_25 & (~ IN2[44]) | select_ne_25 & (~ IN2[45])  );
    wire logic pp_25_46;
    assign pp_25_46 = (select_e_25 & IN2[46] | select_2x_25 & IN2[45] | select_n2x_25 & (~ IN2[45]) | select_ne_25 & (~ IN2[46])  );
    wire logic pp_25_47;
    assign pp_25_47 = (select_e_25 & IN2[47] | select_2x_25 & IN2[46] | select_n2x_25 & (~ IN2[46]) | select_ne_25 & (~ IN2[47])  );
    wire logic pp_25_48;
    assign pp_25_48 = (select_e_25 & IN2[48] | select_2x_25 & IN2[47] | select_n2x_25 & (~ IN2[47]) | select_ne_25 & (~ IN2[48])  );
    wire logic pp_25_49;
    assign pp_25_49 = (select_e_25 & IN2[49] | select_2x_25 & IN2[48] | select_n2x_25 & (~ IN2[48]) | select_ne_25 & (~ IN2[49])  );
    wire logic pp_25_50;
    assign pp_25_50 = (select_e_25 & IN2[50] | select_2x_25 & IN2[49] | select_n2x_25 & (~ IN2[49]) | select_ne_25 & (~ IN2[50])  );
    wire logic pp_25_51;
    assign pp_25_51 = (select_e_25 & IN2[51] | select_2x_25 & IN2[50] | select_n2x_25 & (~ IN2[50]) | select_ne_25 & (~ IN2[51])  );
    wire logic pp_25_52;
    assign pp_25_52 = (select_e_25 & IN2[52] | select_2x_25 & IN2[51] | select_n2x_25 & (~ IN2[51]) | select_ne_25 & (~ IN2[52])  );
    wire logic pp_25_53;
    assign pp_25_53 = (select_e_25 & IN2[53] | select_2x_25 & IN2[52] | select_n2x_25 & (~ IN2[52]) | select_ne_25 & (~ IN2[53])  );
    wire logic pp_25_54;
    assign pp_25_54 = (select_e_25 & IN2[54] | select_2x_25 & IN2[53] | select_n2x_25 & (~ IN2[53]) | select_ne_25 & (~ IN2[54])  );
    wire logic pp_25_55;
    assign pp_25_55 = (select_e_25 & IN2[55] | select_2x_25 & IN2[54] | select_n2x_25 & (~ IN2[54]) | select_ne_25 & (~ IN2[55])  );
    wire logic pp_25_56;
    assign pp_25_56 = (select_e_25 & IN2[56] | select_2x_25 & IN2[55] | select_n2x_25 & (~ IN2[55]) | select_ne_25 & (~ IN2[56])  );
    wire logic pp_25_57;
    assign pp_25_57 = (select_e_25 & IN2[57] | select_2x_25 & IN2[56] | select_n2x_25 & (~ IN2[56]) | select_ne_25 & (~ IN2[57])  );
    wire logic pp_25_58;
    assign pp_25_58 = (select_e_25 & IN2[58] | select_2x_25 & IN2[57] | select_n2x_25 & (~ IN2[57]) | select_ne_25 & (~ IN2[58])  );
    wire logic pp_25_59;
    assign pp_25_59 = (select_e_25 & IN2[59] | select_2x_25 & IN2[58] | select_n2x_25 & (~ IN2[58]) | select_ne_25 & (~ IN2[59])  );
    wire logic pp_25_60;
    assign pp_25_60 = (select_e_25 & IN2[60] | select_2x_25 & IN2[59] | select_n2x_25 & (~ IN2[59]) | select_ne_25 & (~ IN2[60])  );
    wire logic pp_25_61;
    assign pp_25_61 = (select_e_25 & IN2[61] | select_2x_25 & IN2[60] | select_n2x_25 & (~ IN2[60]) | select_ne_25 & (~ IN2[61])  );
    wire logic pp_25_62;
    assign pp_25_62 = (select_e_25 & IN2[62] | select_2x_25 & IN2[61] | select_n2x_25 & (~ IN2[61]) | select_ne_25 & (~ IN2[62])  );
    wire logic pp_25_63;
    assign pp_25_63 = (select_e_25 & IN2[63] | select_2x_25 & IN2[62] | select_n2x_25 & (~ IN2[62]) | select_ne_25 & (~ IN2[63])  );
    wire logic pp_25_64;
    assign pp_25_64 = (select_e_25 & IN2[63] | select_2x_25 & IN2[63] | select_n2x_25 & (~ IN2[63]) | select_ne_25 & (~ IN2[63])  );
    wire logic pp_25_65;
    assign pp_25_65 = ~ (select_e_25 & IN2[63] | select_2x_25 & IN2[63] | select_n2x_25 & (~ IN2[63]) | select_ne_25 & (~ IN2[63])  );
    assign tcomp25 = select_ne_25 | select_n2x_25;
    
    // Signed Booth Radix-4 Partial Products Row 27
    wire logic select_e_26, select_ne_26, select_2x_26, tcomp26, select_n2x_26;
    assign select_e_26 = ((~ IN1[53]) & (IN1[52] ^ IN1[51]));
    assign select_ne_26 = IN1[53] &  (IN1[52] ^ IN1[51]);
    assign select_2x_26 = (~ IN1[53]) & IN1[52] & IN1[51];
    assign select_n2x_26 = IN1[53] & (~ IN1[52]) & (~ IN1[51]);
    wire logic pp_26_0;
    assign pp_26_0 = (select_e_26 & IN2[0] | select_2x_26 & 1'b0 | select_n2x_26 & 1'b1 | select_ne_26 & (~ IN2[0])  );
    wire logic pp_26_1;
    assign pp_26_1 = (select_e_26 & IN2[1] | select_2x_26 & IN2[0] | select_n2x_26 & (~ IN2[0]) | select_ne_26 & (~ IN2[1])  );
    wire logic pp_26_2;
    assign pp_26_2 = (select_e_26 & IN2[2] | select_2x_26 & IN2[1] | select_n2x_26 & (~ IN2[1]) | select_ne_26 & (~ IN2[2])  );
    wire logic pp_26_3;
    assign pp_26_3 = (select_e_26 & IN2[3] | select_2x_26 & IN2[2] | select_n2x_26 & (~ IN2[2]) | select_ne_26 & (~ IN2[3])  );
    wire logic pp_26_4;
    assign pp_26_4 = (select_e_26 & IN2[4] | select_2x_26 & IN2[3] | select_n2x_26 & (~ IN2[3]) | select_ne_26 & (~ IN2[4])  );
    wire logic pp_26_5;
    assign pp_26_5 = (select_e_26 & IN2[5] | select_2x_26 & IN2[4] | select_n2x_26 & (~ IN2[4]) | select_ne_26 & (~ IN2[5])  );
    wire logic pp_26_6;
    assign pp_26_6 = (select_e_26 & IN2[6] | select_2x_26 & IN2[5] | select_n2x_26 & (~ IN2[5]) | select_ne_26 & (~ IN2[6])  );
    wire logic pp_26_7;
    assign pp_26_7 = (select_e_26 & IN2[7] | select_2x_26 & IN2[6] | select_n2x_26 & (~ IN2[6]) | select_ne_26 & (~ IN2[7])  );
    wire logic pp_26_8;
    assign pp_26_8 = (select_e_26 & IN2[8] | select_2x_26 & IN2[7] | select_n2x_26 & (~ IN2[7]) | select_ne_26 & (~ IN2[8])  );
    wire logic pp_26_9;
    assign pp_26_9 = (select_e_26 & IN2[9] | select_2x_26 & IN2[8] | select_n2x_26 & (~ IN2[8]) | select_ne_26 & (~ IN2[9])  );
    wire logic pp_26_10;
    assign pp_26_10 = (select_e_26 & IN2[10] | select_2x_26 & IN2[9] | select_n2x_26 & (~ IN2[9]) | select_ne_26 & (~ IN2[10])  );
    wire logic pp_26_11;
    assign pp_26_11 = (select_e_26 & IN2[11] | select_2x_26 & IN2[10] | select_n2x_26 & (~ IN2[10]) | select_ne_26 & (~ IN2[11])  );
    wire logic pp_26_12;
    assign pp_26_12 = (select_e_26 & IN2[12] | select_2x_26 & IN2[11] | select_n2x_26 & (~ IN2[11]) | select_ne_26 & (~ IN2[12])  );
    wire logic pp_26_13;
    assign pp_26_13 = (select_e_26 & IN2[13] | select_2x_26 & IN2[12] | select_n2x_26 & (~ IN2[12]) | select_ne_26 & (~ IN2[13])  );
    wire logic pp_26_14;
    assign pp_26_14 = (select_e_26 & IN2[14] | select_2x_26 & IN2[13] | select_n2x_26 & (~ IN2[13]) | select_ne_26 & (~ IN2[14])  );
    wire logic pp_26_15;
    assign pp_26_15 = (select_e_26 & IN2[15] | select_2x_26 & IN2[14] | select_n2x_26 & (~ IN2[14]) | select_ne_26 & (~ IN2[15])  );
    wire logic pp_26_16;
    assign pp_26_16 = (select_e_26 & IN2[16] | select_2x_26 & IN2[15] | select_n2x_26 & (~ IN2[15]) | select_ne_26 & (~ IN2[16])  );
    wire logic pp_26_17;
    assign pp_26_17 = (select_e_26 & IN2[17] | select_2x_26 & IN2[16] | select_n2x_26 & (~ IN2[16]) | select_ne_26 & (~ IN2[17])  );
    wire logic pp_26_18;
    assign pp_26_18 = (select_e_26 & IN2[18] | select_2x_26 & IN2[17] | select_n2x_26 & (~ IN2[17]) | select_ne_26 & (~ IN2[18])  );
    wire logic pp_26_19;
    assign pp_26_19 = (select_e_26 & IN2[19] | select_2x_26 & IN2[18] | select_n2x_26 & (~ IN2[18]) | select_ne_26 & (~ IN2[19])  );
    wire logic pp_26_20;
    assign pp_26_20 = (select_e_26 & IN2[20] | select_2x_26 & IN2[19] | select_n2x_26 & (~ IN2[19]) | select_ne_26 & (~ IN2[20])  );
    wire logic pp_26_21;
    assign pp_26_21 = (select_e_26 & IN2[21] | select_2x_26 & IN2[20] | select_n2x_26 & (~ IN2[20]) | select_ne_26 & (~ IN2[21])  );
    wire logic pp_26_22;
    assign pp_26_22 = (select_e_26 & IN2[22] | select_2x_26 & IN2[21] | select_n2x_26 & (~ IN2[21]) | select_ne_26 & (~ IN2[22])  );
    wire logic pp_26_23;
    assign pp_26_23 = (select_e_26 & IN2[23] | select_2x_26 & IN2[22] | select_n2x_26 & (~ IN2[22]) | select_ne_26 & (~ IN2[23])  );
    wire logic pp_26_24;
    assign pp_26_24 = (select_e_26 & IN2[24] | select_2x_26 & IN2[23] | select_n2x_26 & (~ IN2[23]) | select_ne_26 & (~ IN2[24])  );
    wire logic pp_26_25;
    assign pp_26_25 = (select_e_26 & IN2[25] | select_2x_26 & IN2[24] | select_n2x_26 & (~ IN2[24]) | select_ne_26 & (~ IN2[25])  );
    wire logic pp_26_26;
    assign pp_26_26 = (select_e_26 & IN2[26] | select_2x_26 & IN2[25] | select_n2x_26 & (~ IN2[25]) | select_ne_26 & (~ IN2[26])  );
    wire logic pp_26_27;
    assign pp_26_27 = (select_e_26 & IN2[27] | select_2x_26 & IN2[26] | select_n2x_26 & (~ IN2[26]) | select_ne_26 & (~ IN2[27])  );
    wire logic pp_26_28;
    assign pp_26_28 = (select_e_26 & IN2[28] | select_2x_26 & IN2[27] | select_n2x_26 & (~ IN2[27]) | select_ne_26 & (~ IN2[28])  );
    wire logic pp_26_29;
    assign pp_26_29 = (select_e_26 & IN2[29] | select_2x_26 & IN2[28] | select_n2x_26 & (~ IN2[28]) | select_ne_26 & (~ IN2[29])  );
    wire logic pp_26_30;
    assign pp_26_30 = (select_e_26 & IN2[30] | select_2x_26 & IN2[29] | select_n2x_26 & (~ IN2[29]) | select_ne_26 & (~ IN2[30])  );
    wire logic pp_26_31;
    assign pp_26_31 = (select_e_26 & IN2[31] | select_2x_26 & IN2[30] | select_n2x_26 & (~ IN2[30]) | select_ne_26 & (~ IN2[31])  );
    wire logic pp_26_32;
    assign pp_26_32 = (select_e_26 & IN2[32] | select_2x_26 & IN2[31] | select_n2x_26 & (~ IN2[31]) | select_ne_26 & (~ IN2[32])  );
    wire logic pp_26_33;
    assign pp_26_33 = (select_e_26 & IN2[33] | select_2x_26 & IN2[32] | select_n2x_26 & (~ IN2[32]) | select_ne_26 & (~ IN2[33])  );
    wire logic pp_26_34;
    assign pp_26_34 = (select_e_26 & IN2[34] | select_2x_26 & IN2[33] | select_n2x_26 & (~ IN2[33]) | select_ne_26 & (~ IN2[34])  );
    wire logic pp_26_35;
    assign pp_26_35 = (select_e_26 & IN2[35] | select_2x_26 & IN2[34] | select_n2x_26 & (~ IN2[34]) | select_ne_26 & (~ IN2[35])  );
    wire logic pp_26_36;
    assign pp_26_36 = (select_e_26 & IN2[36] | select_2x_26 & IN2[35] | select_n2x_26 & (~ IN2[35]) | select_ne_26 & (~ IN2[36])  );
    wire logic pp_26_37;
    assign pp_26_37 = (select_e_26 & IN2[37] | select_2x_26 & IN2[36] | select_n2x_26 & (~ IN2[36]) | select_ne_26 & (~ IN2[37])  );
    wire logic pp_26_38;
    assign pp_26_38 = (select_e_26 & IN2[38] | select_2x_26 & IN2[37] | select_n2x_26 & (~ IN2[37]) | select_ne_26 & (~ IN2[38])  );
    wire logic pp_26_39;
    assign pp_26_39 = (select_e_26 & IN2[39] | select_2x_26 & IN2[38] | select_n2x_26 & (~ IN2[38]) | select_ne_26 & (~ IN2[39])  );
    wire logic pp_26_40;
    assign pp_26_40 = (select_e_26 & IN2[40] | select_2x_26 & IN2[39] | select_n2x_26 & (~ IN2[39]) | select_ne_26 & (~ IN2[40])  );
    wire logic pp_26_41;
    assign pp_26_41 = (select_e_26 & IN2[41] | select_2x_26 & IN2[40] | select_n2x_26 & (~ IN2[40]) | select_ne_26 & (~ IN2[41])  );
    wire logic pp_26_42;
    assign pp_26_42 = (select_e_26 & IN2[42] | select_2x_26 & IN2[41] | select_n2x_26 & (~ IN2[41]) | select_ne_26 & (~ IN2[42])  );
    wire logic pp_26_43;
    assign pp_26_43 = (select_e_26 & IN2[43] | select_2x_26 & IN2[42] | select_n2x_26 & (~ IN2[42]) | select_ne_26 & (~ IN2[43])  );
    wire logic pp_26_44;
    assign pp_26_44 = (select_e_26 & IN2[44] | select_2x_26 & IN2[43] | select_n2x_26 & (~ IN2[43]) | select_ne_26 & (~ IN2[44])  );
    wire logic pp_26_45;
    assign pp_26_45 = (select_e_26 & IN2[45] | select_2x_26 & IN2[44] | select_n2x_26 & (~ IN2[44]) | select_ne_26 & (~ IN2[45])  );
    wire logic pp_26_46;
    assign pp_26_46 = (select_e_26 & IN2[46] | select_2x_26 & IN2[45] | select_n2x_26 & (~ IN2[45]) | select_ne_26 & (~ IN2[46])  );
    wire logic pp_26_47;
    assign pp_26_47 = (select_e_26 & IN2[47] | select_2x_26 & IN2[46] | select_n2x_26 & (~ IN2[46]) | select_ne_26 & (~ IN2[47])  );
    wire logic pp_26_48;
    assign pp_26_48 = (select_e_26 & IN2[48] | select_2x_26 & IN2[47] | select_n2x_26 & (~ IN2[47]) | select_ne_26 & (~ IN2[48])  );
    wire logic pp_26_49;
    assign pp_26_49 = (select_e_26 & IN2[49] | select_2x_26 & IN2[48] | select_n2x_26 & (~ IN2[48]) | select_ne_26 & (~ IN2[49])  );
    wire logic pp_26_50;
    assign pp_26_50 = (select_e_26 & IN2[50] | select_2x_26 & IN2[49] | select_n2x_26 & (~ IN2[49]) | select_ne_26 & (~ IN2[50])  );
    wire logic pp_26_51;
    assign pp_26_51 = (select_e_26 & IN2[51] | select_2x_26 & IN2[50] | select_n2x_26 & (~ IN2[50]) | select_ne_26 & (~ IN2[51])  );
    wire logic pp_26_52;
    assign pp_26_52 = (select_e_26 & IN2[52] | select_2x_26 & IN2[51] | select_n2x_26 & (~ IN2[51]) | select_ne_26 & (~ IN2[52])  );
    wire logic pp_26_53;
    assign pp_26_53 = (select_e_26 & IN2[53] | select_2x_26 & IN2[52] | select_n2x_26 & (~ IN2[52]) | select_ne_26 & (~ IN2[53])  );
    wire logic pp_26_54;
    assign pp_26_54 = (select_e_26 & IN2[54] | select_2x_26 & IN2[53] | select_n2x_26 & (~ IN2[53]) | select_ne_26 & (~ IN2[54])  );
    wire logic pp_26_55;
    assign pp_26_55 = (select_e_26 & IN2[55] | select_2x_26 & IN2[54] | select_n2x_26 & (~ IN2[54]) | select_ne_26 & (~ IN2[55])  );
    wire logic pp_26_56;
    assign pp_26_56 = (select_e_26 & IN2[56] | select_2x_26 & IN2[55] | select_n2x_26 & (~ IN2[55]) | select_ne_26 & (~ IN2[56])  );
    wire logic pp_26_57;
    assign pp_26_57 = (select_e_26 & IN2[57] | select_2x_26 & IN2[56] | select_n2x_26 & (~ IN2[56]) | select_ne_26 & (~ IN2[57])  );
    wire logic pp_26_58;
    assign pp_26_58 = (select_e_26 & IN2[58] | select_2x_26 & IN2[57] | select_n2x_26 & (~ IN2[57]) | select_ne_26 & (~ IN2[58])  );
    wire logic pp_26_59;
    assign pp_26_59 = (select_e_26 & IN2[59] | select_2x_26 & IN2[58] | select_n2x_26 & (~ IN2[58]) | select_ne_26 & (~ IN2[59])  );
    wire logic pp_26_60;
    assign pp_26_60 = (select_e_26 & IN2[60] | select_2x_26 & IN2[59] | select_n2x_26 & (~ IN2[59]) | select_ne_26 & (~ IN2[60])  );
    wire logic pp_26_61;
    assign pp_26_61 = (select_e_26 & IN2[61] | select_2x_26 & IN2[60] | select_n2x_26 & (~ IN2[60]) | select_ne_26 & (~ IN2[61])  );
    wire logic pp_26_62;
    assign pp_26_62 = (select_e_26 & IN2[62] | select_2x_26 & IN2[61] | select_n2x_26 & (~ IN2[61]) | select_ne_26 & (~ IN2[62])  );
    wire logic pp_26_63;
    assign pp_26_63 = (select_e_26 & IN2[63] | select_2x_26 & IN2[62] | select_n2x_26 & (~ IN2[62]) | select_ne_26 & (~ IN2[63])  );
    wire logic pp_26_64;
    assign pp_26_64 = (select_e_26 & IN2[63] | select_2x_26 & IN2[63] | select_n2x_26 & (~ IN2[63]) | select_ne_26 & (~ IN2[63])  );
    wire logic pp_26_65;
    assign pp_26_65 = ~ (select_e_26 & IN2[63] | select_2x_26 & IN2[63] | select_n2x_26 & (~ IN2[63]) | select_ne_26 & (~ IN2[63])  );
    assign tcomp26 = select_ne_26 | select_n2x_26;
    
    // Signed Booth Radix-4 Partial Products Row 28
    wire logic select_e_27, select_ne_27, select_2x_27, tcomp27, select_n2x_27;
    assign select_e_27 = ((~ IN1[55]) & (IN1[54] ^ IN1[53]));
    assign select_ne_27 = IN1[55] &  (IN1[54] ^ IN1[53]);
    assign select_2x_27 = (~ IN1[55]) & IN1[54] & IN1[53];
    assign select_n2x_27 = IN1[55] & (~ IN1[54]) & (~ IN1[53]);
    wire logic pp_27_0;
    assign pp_27_0 = (select_e_27 & IN2[0] | select_2x_27 & 1'b0 | select_n2x_27 & 1'b1 | select_ne_27 & (~ IN2[0])  );
    wire logic pp_27_1;
    assign pp_27_1 = (select_e_27 & IN2[1] | select_2x_27 & IN2[0] | select_n2x_27 & (~ IN2[0]) | select_ne_27 & (~ IN2[1])  );
    wire logic pp_27_2;
    assign pp_27_2 = (select_e_27 & IN2[2] | select_2x_27 & IN2[1] | select_n2x_27 & (~ IN2[1]) | select_ne_27 & (~ IN2[2])  );
    wire logic pp_27_3;
    assign pp_27_3 = (select_e_27 & IN2[3] | select_2x_27 & IN2[2] | select_n2x_27 & (~ IN2[2]) | select_ne_27 & (~ IN2[3])  );
    wire logic pp_27_4;
    assign pp_27_4 = (select_e_27 & IN2[4] | select_2x_27 & IN2[3] | select_n2x_27 & (~ IN2[3]) | select_ne_27 & (~ IN2[4])  );
    wire logic pp_27_5;
    assign pp_27_5 = (select_e_27 & IN2[5] | select_2x_27 & IN2[4] | select_n2x_27 & (~ IN2[4]) | select_ne_27 & (~ IN2[5])  );
    wire logic pp_27_6;
    assign pp_27_6 = (select_e_27 & IN2[6] | select_2x_27 & IN2[5] | select_n2x_27 & (~ IN2[5]) | select_ne_27 & (~ IN2[6])  );
    wire logic pp_27_7;
    assign pp_27_7 = (select_e_27 & IN2[7] | select_2x_27 & IN2[6] | select_n2x_27 & (~ IN2[6]) | select_ne_27 & (~ IN2[7])  );
    wire logic pp_27_8;
    assign pp_27_8 = (select_e_27 & IN2[8] | select_2x_27 & IN2[7] | select_n2x_27 & (~ IN2[7]) | select_ne_27 & (~ IN2[8])  );
    wire logic pp_27_9;
    assign pp_27_9 = (select_e_27 & IN2[9] | select_2x_27 & IN2[8] | select_n2x_27 & (~ IN2[8]) | select_ne_27 & (~ IN2[9])  );
    wire logic pp_27_10;
    assign pp_27_10 = (select_e_27 & IN2[10] | select_2x_27 & IN2[9] | select_n2x_27 & (~ IN2[9]) | select_ne_27 & (~ IN2[10])  );
    wire logic pp_27_11;
    assign pp_27_11 = (select_e_27 & IN2[11] | select_2x_27 & IN2[10] | select_n2x_27 & (~ IN2[10]) | select_ne_27 & (~ IN2[11])  );
    wire logic pp_27_12;
    assign pp_27_12 = (select_e_27 & IN2[12] | select_2x_27 & IN2[11] | select_n2x_27 & (~ IN2[11]) | select_ne_27 & (~ IN2[12])  );
    wire logic pp_27_13;
    assign pp_27_13 = (select_e_27 & IN2[13] | select_2x_27 & IN2[12] | select_n2x_27 & (~ IN2[12]) | select_ne_27 & (~ IN2[13])  );
    wire logic pp_27_14;
    assign pp_27_14 = (select_e_27 & IN2[14] | select_2x_27 & IN2[13] | select_n2x_27 & (~ IN2[13]) | select_ne_27 & (~ IN2[14])  );
    wire logic pp_27_15;
    assign pp_27_15 = (select_e_27 & IN2[15] | select_2x_27 & IN2[14] | select_n2x_27 & (~ IN2[14]) | select_ne_27 & (~ IN2[15])  );
    wire logic pp_27_16;
    assign pp_27_16 = (select_e_27 & IN2[16] | select_2x_27 & IN2[15] | select_n2x_27 & (~ IN2[15]) | select_ne_27 & (~ IN2[16])  );
    wire logic pp_27_17;
    assign pp_27_17 = (select_e_27 & IN2[17] | select_2x_27 & IN2[16] | select_n2x_27 & (~ IN2[16]) | select_ne_27 & (~ IN2[17])  );
    wire logic pp_27_18;
    assign pp_27_18 = (select_e_27 & IN2[18] | select_2x_27 & IN2[17] | select_n2x_27 & (~ IN2[17]) | select_ne_27 & (~ IN2[18])  );
    wire logic pp_27_19;
    assign pp_27_19 = (select_e_27 & IN2[19] | select_2x_27 & IN2[18] | select_n2x_27 & (~ IN2[18]) | select_ne_27 & (~ IN2[19])  );
    wire logic pp_27_20;
    assign pp_27_20 = (select_e_27 & IN2[20] | select_2x_27 & IN2[19] | select_n2x_27 & (~ IN2[19]) | select_ne_27 & (~ IN2[20])  );
    wire logic pp_27_21;
    assign pp_27_21 = (select_e_27 & IN2[21] | select_2x_27 & IN2[20] | select_n2x_27 & (~ IN2[20]) | select_ne_27 & (~ IN2[21])  );
    wire logic pp_27_22;
    assign pp_27_22 = (select_e_27 & IN2[22] | select_2x_27 & IN2[21] | select_n2x_27 & (~ IN2[21]) | select_ne_27 & (~ IN2[22])  );
    wire logic pp_27_23;
    assign pp_27_23 = (select_e_27 & IN2[23] | select_2x_27 & IN2[22] | select_n2x_27 & (~ IN2[22]) | select_ne_27 & (~ IN2[23])  );
    wire logic pp_27_24;
    assign pp_27_24 = (select_e_27 & IN2[24] | select_2x_27 & IN2[23] | select_n2x_27 & (~ IN2[23]) | select_ne_27 & (~ IN2[24])  );
    wire logic pp_27_25;
    assign pp_27_25 = (select_e_27 & IN2[25] | select_2x_27 & IN2[24] | select_n2x_27 & (~ IN2[24]) | select_ne_27 & (~ IN2[25])  );
    wire logic pp_27_26;
    assign pp_27_26 = (select_e_27 & IN2[26] | select_2x_27 & IN2[25] | select_n2x_27 & (~ IN2[25]) | select_ne_27 & (~ IN2[26])  );
    wire logic pp_27_27;
    assign pp_27_27 = (select_e_27 & IN2[27] | select_2x_27 & IN2[26] | select_n2x_27 & (~ IN2[26]) | select_ne_27 & (~ IN2[27])  );
    wire logic pp_27_28;
    assign pp_27_28 = (select_e_27 & IN2[28] | select_2x_27 & IN2[27] | select_n2x_27 & (~ IN2[27]) | select_ne_27 & (~ IN2[28])  );
    wire logic pp_27_29;
    assign pp_27_29 = (select_e_27 & IN2[29] | select_2x_27 & IN2[28] | select_n2x_27 & (~ IN2[28]) | select_ne_27 & (~ IN2[29])  );
    wire logic pp_27_30;
    assign pp_27_30 = (select_e_27 & IN2[30] | select_2x_27 & IN2[29] | select_n2x_27 & (~ IN2[29]) | select_ne_27 & (~ IN2[30])  );
    wire logic pp_27_31;
    assign pp_27_31 = (select_e_27 & IN2[31] | select_2x_27 & IN2[30] | select_n2x_27 & (~ IN2[30]) | select_ne_27 & (~ IN2[31])  );
    wire logic pp_27_32;
    assign pp_27_32 = (select_e_27 & IN2[32] | select_2x_27 & IN2[31] | select_n2x_27 & (~ IN2[31]) | select_ne_27 & (~ IN2[32])  );
    wire logic pp_27_33;
    assign pp_27_33 = (select_e_27 & IN2[33] | select_2x_27 & IN2[32] | select_n2x_27 & (~ IN2[32]) | select_ne_27 & (~ IN2[33])  );
    wire logic pp_27_34;
    assign pp_27_34 = (select_e_27 & IN2[34] | select_2x_27 & IN2[33] | select_n2x_27 & (~ IN2[33]) | select_ne_27 & (~ IN2[34])  );
    wire logic pp_27_35;
    assign pp_27_35 = (select_e_27 & IN2[35] | select_2x_27 & IN2[34] | select_n2x_27 & (~ IN2[34]) | select_ne_27 & (~ IN2[35])  );
    wire logic pp_27_36;
    assign pp_27_36 = (select_e_27 & IN2[36] | select_2x_27 & IN2[35] | select_n2x_27 & (~ IN2[35]) | select_ne_27 & (~ IN2[36])  );
    wire logic pp_27_37;
    assign pp_27_37 = (select_e_27 & IN2[37] | select_2x_27 & IN2[36] | select_n2x_27 & (~ IN2[36]) | select_ne_27 & (~ IN2[37])  );
    wire logic pp_27_38;
    assign pp_27_38 = (select_e_27 & IN2[38] | select_2x_27 & IN2[37] | select_n2x_27 & (~ IN2[37]) | select_ne_27 & (~ IN2[38])  );
    wire logic pp_27_39;
    assign pp_27_39 = (select_e_27 & IN2[39] | select_2x_27 & IN2[38] | select_n2x_27 & (~ IN2[38]) | select_ne_27 & (~ IN2[39])  );
    wire logic pp_27_40;
    assign pp_27_40 = (select_e_27 & IN2[40] | select_2x_27 & IN2[39] | select_n2x_27 & (~ IN2[39]) | select_ne_27 & (~ IN2[40])  );
    wire logic pp_27_41;
    assign pp_27_41 = (select_e_27 & IN2[41] | select_2x_27 & IN2[40] | select_n2x_27 & (~ IN2[40]) | select_ne_27 & (~ IN2[41])  );
    wire logic pp_27_42;
    assign pp_27_42 = (select_e_27 & IN2[42] | select_2x_27 & IN2[41] | select_n2x_27 & (~ IN2[41]) | select_ne_27 & (~ IN2[42])  );
    wire logic pp_27_43;
    assign pp_27_43 = (select_e_27 & IN2[43] | select_2x_27 & IN2[42] | select_n2x_27 & (~ IN2[42]) | select_ne_27 & (~ IN2[43])  );
    wire logic pp_27_44;
    assign pp_27_44 = (select_e_27 & IN2[44] | select_2x_27 & IN2[43] | select_n2x_27 & (~ IN2[43]) | select_ne_27 & (~ IN2[44])  );
    wire logic pp_27_45;
    assign pp_27_45 = (select_e_27 & IN2[45] | select_2x_27 & IN2[44] | select_n2x_27 & (~ IN2[44]) | select_ne_27 & (~ IN2[45])  );
    wire logic pp_27_46;
    assign pp_27_46 = (select_e_27 & IN2[46] | select_2x_27 & IN2[45] | select_n2x_27 & (~ IN2[45]) | select_ne_27 & (~ IN2[46])  );
    wire logic pp_27_47;
    assign pp_27_47 = (select_e_27 & IN2[47] | select_2x_27 & IN2[46] | select_n2x_27 & (~ IN2[46]) | select_ne_27 & (~ IN2[47])  );
    wire logic pp_27_48;
    assign pp_27_48 = (select_e_27 & IN2[48] | select_2x_27 & IN2[47] | select_n2x_27 & (~ IN2[47]) | select_ne_27 & (~ IN2[48])  );
    wire logic pp_27_49;
    assign pp_27_49 = (select_e_27 & IN2[49] | select_2x_27 & IN2[48] | select_n2x_27 & (~ IN2[48]) | select_ne_27 & (~ IN2[49])  );
    wire logic pp_27_50;
    assign pp_27_50 = (select_e_27 & IN2[50] | select_2x_27 & IN2[49] | select_n2x_27 & (~ IN2[49]) | select_ne_27 & (~ IN2[50])  );
    wire logic pp_27_51;
    assign pp_27_51 = (select_e_27 & IN2[51] | select_2x_27 & IN2[50] | select_n2x_27 & (~ IN2[50]) | select_ne_27 & (~ IN2[51])  );
    wire logic pp_27_52;
    assign pp_27_52 = (select_e_27 & IN2[52] | select_2x_27 & IN2[51] | select_n2x_27 & (~ IN2[51]) | select_ne_27 & (~ IN2[52])  );
    wire logic pp_27_53;
    assign pp_27_53 = (select_e_27 & IN2[53] | select_2x_27 & IN2[52] | select_n2x_27 & (~ IN2[52]) | select_ne_27 & (~ IN2[53])  );
    wire logic pp_27_54;
    assign pp_27_54 = (select_e_27 & IN2[54] | select_2x_27 & IN2[53] | select_n2x_27 & (~ IN2[53]) | select_ne_27 & (~ IN2[54])  );
    wire logic pp_27_55;
    assign pp_27_55 = (select_e_27 & IN2[55] | select_2x_27 & IN2[54] | select_n2x_27 & (~ IN2[54]) | select_ne_27 & (~ IN2[55])  );
    wire logic pp_27_56;
    assign pp_27_56 = (select_e_27 & IN2[56] | select_2x_27 & IN2[55] | select_n2x_27 & (~ IN2[55]) | select_ne_27 & (~ IN2[56])  );
    wire logic pp_27_57;
    assign pp_27_57 = (select_e_27 & IN2[57] | select_2x_27 & IN2[56] | select_n2x_27 & (~ IN2[56]) | select_ne_27 & (~ IN2[57])  );
    wire logic pp_27_58;
    assign pp_27_58 = (select_e_27 & IN2[58] | select_2x_27 & IN2[57] | select_n2x_27 & (~ IN2[57]) | select_ne_27 & (~ IN2[58])  );
    wire logic pp_27_59;
    assign pp_27_59 = (select_e_27 & IN2[59] | select_2x_27 & IN2[58] | select_n2x_27 & (~ IN2[58]) | select_ne_27 & (~ IN2[59])  );
    wire logic pp_27_60;
    assign pp_27_60 = (select_e_27 & IN2[60] | select_2x_27 & IN2[59] | select_n2x_27 & (~ IN2[59]) | select_ne_27 & (~ IN2[60])  );
    wire logic pp_27_61;
    assign pp_27_61 = (select_e_27 & IN2[61] | select_2x_27 & IN2[60] | select_n2x_27 & (~ IN2[60]) | select_ne_27 & (~ IN2[61])  );
    wire logic pp_27_62;
    assign pp_27_62 = (select_e_27 & IN2[62] | select_2x_27 & IN2[61] | select_n2x_27 & (~ IN2[61]) | select_ne_27 & (~ IN2[62])  );
    wire logic pp_27_63;
    assign pp_27_63 = (select_e_27 & IN2[63] | select_2x_27 & IN2[62] | select_n2x_27 & (~ IN2[62]) | select_ne_27 & (~ IN2[63])  );
    wire logic pp_27_64;
    assign pp_27_64 = (select_e_27 & IN2[63] | select_2x_27 & IN2[63] | select_n2x_27 & (~ IN2[63]) | select_ne_27 & (~ IN2[63])  );
    wire logic pp_27_65;
    assign pp_27_65 = ~ (select_e_27 & IN2[63] | select_2x_27 & IN2[63] | select_n2x_27 & (~ IN2[63]) | select_ne_27 & (~ IN2[63])  );
    assign tcomp27 = select_ne_27 | select_n2x_27;
    
    // Signed Booth Radix-4 Partial Products Row 29
    wire logic select_e_28, select_ne_28, select_2x_28, tcomp28, select_n2x_28;
    assign select_e_28 = ((~ IN1[57]) & (IN1[56] ^ IN1[55]));
    assign select_ne_28 = IN1[57] &  (IN1[56] ^ IN1[55]);
    assign select_2x_28 = (~ IN1[57]) & IN1[56] & IN1[55];
    assign select_n2x_28 = IN1[57] & (~ IN1[56]) & (~ IN1[55]);
    wire logic pp_28_0;
    assign pp_28_0 = (select_e_28 & IN2[0] | select_2x_28 & 1'b0 | select_n2x_28 & 1'b1 | select_ne_28 & (~ IN2[0])  );
    wire logic pp_28_1;
    assign pp_28_1 = (select_e_28 & IN2[1] | select_2x_28 & IN2[0] | select_n2x_28 & (~ IN2[0]) | select_ne_28 & (~ IN2[1])  );
    wire logic pp_28_2;
    assign pp_28_2 = (select_e_28 & IN2[2] | select_2x_28 & IN2[1] | select_n2x_28 & (~ IN2[1]) | select_ne_28 & (~ IN2[2])  );
    wire logic pp_28_3;
    assign pp_28_3 = (select_e_28 & IN2[3] | select_2x_28 & IN2[2] | select_n2x_28 & (~ IN2[2]) | select_ne_28 & (~ IN2[3])  );
    wire logic pp_28_4;
    assign pp_28_4 = (select_e_28 & IN2[4] | select_2x_28 & IN2[3] | select_n2x_28 & (~ IN2[3]) | select_ne_28 & (~ IN2[4])  );
    wire logic pp_28_5;
    assign pp_28_5 = (select_e_28 & IN2[5] | select_2x_28 & IN2[4] | select_n2x_28 & (~ IN2[4]) | select_ne_28 & (~ IN2[5])  );
    wire logic pp_28_6;
    assign pp_28_6 = (select_e_28 & IN2[6] | select_2x_28 & IN2[5] | select_n2x_28 & (~ IN2[5]) | select_ne_28 & (~ IN2[6])  );
    wire logic pp_28_7;
    assign pp_28_7 = (select_e_28 & IN2[7] | select_2x_28 & IN2[6] | select_n2x_28 & (~ IN2[6]) | select_ne_28 & (~ IN2[7])  );
    wire logic pp_28_8;
    assign pp_28_8 = (select_e_28 & IN2[8] | select_2x_28 & IN2[7] | select_n2x_28 & (~ IN2[7]) | select_ne_28 & (~ IN2[8])  );
    wire logic pp_28_9;
    assign pp_28_9 = (select_e_28 & IN2[9] | select_2x_28 & IN2[8] | select_n2x_28 & (~ IN2[8]) | select_ne_28 & (~ IN2[9])  );
    wire logic pp_28_10;
    assign pp_28_10 = (select_e_28 & IN2[10] | select_2x_28 & IN2[9] | select_n2x_28 & (~ IN2[9]) | select_ne_28 & (~ IN2[10])  );
    wire logic pp_28_11;
    assign pp_28_11 = (select_e_28 & IN2[11] | select_2x_28 & IN2[10] | select_n2x_28 & (~ IN2[10]) | select_ne_28 & (~ IN2[11])  );
    wire logic pp_28_12;
    assign pp_28_12 = (select_e_28 & IN2[12] | select_2x_28 & IN2[11] | select_n2x_28 & (~ IN2[11]) | select_ne_28 & (~ IN2[12])  );
    wire logic pp_28_13;
    assign pp_28_13 = (select_e_28 & IN2[13] | select_2x_28 & IN2[12] | select_n2x_28 & (~ IN2[12]) | select_ne_28 & (~ IN2[13])  );
    wire logic pp_28_14;
    assign pp_28_14 = (select_e_28 & IN2[14] | select_2x_28 & IN2[13] | select_n2x_28 & (~ IN2[13]) | select_ne_28 & (~ IN2[14])  );
    wire logic pp_28_15;
    assign pp_28_15 = (select_e_28 & IN2[15] | select_2x_28 & IN2[14] | select_n2x_28 & (~ IN2[14]) | select_ne_28 & (~ IN2[15])  );
    wire logic pp_28_16;
    assign pp_28_16 = (select_e_28 & IN2[16] | select_2x_28 & IN2[15] | select_n2x_28 & (~ IN2[15]) | select_ne_28 & (~ IN2[16])  );
    wire logic pp_28_17;
    assign pp_28_17 = (select_e_28 & IN2[17] | select_2x_28 & IN2[16] | select_n2x_28 & (~ IN2[16]) | select_ne_28 & (~ IN2[17])  );
    wire logic pp_28_18;
    assign pp_28_18 = (select_e_28 & IN2[18] | select_2x_28 & IN2[17] | select_n2x_28 & (~ IN2[17]) | select_ne_28 & (~ IN2[18])  );
    wire logic pp_28_19;
    assign pp_28_19 = (select_e_28 & IN2[19] | select_2x_28 & IN2[18] | select_n2x_28 & (~ IN2[18]) | select_ne_28 & (~ IN2[19])  );
    wire logic pp_28_20;
    assign pp_28_20 = (select_e_28 & IN2[20] | select_2x_28 & IN2[19] | select_n2x_28 & (~ IN2[19]) | select_ne_28 & (~ IN2[20])  );
    wire logic pp_28_21;
    assign pp_28_21 = (select_e_28 & IN2[21] | select_2x_28 & IN2[20] | select_n2x_28 & (~ IN2[20]) | select_ne_28 & (~ IN2[21])  );
    wire logic pp_28_22;
    assign pp_28_22 = (select_e_28 & IN2[22] | select_2x_28 & IN2[21] | select_n2x_28 & (~ IN2[21]) | select_ne_28 & (~ IN2[22])  );
    wire logic pp_28_23;
    assign pp_28_23 = (select_e_28 & IN2[23] | select_2x_28 & IN2[22] | select_n2x_28 & (~ IN2[22]) | select_ne_28 & (~ IN2[23])  );
    wire logic pp_28_24;
    assign pp_28_24 = (select_e_28 & IN2[24] | select_2x_28 & IN2[23] | select_n2x_28 & (~ IN2[23]) | select_ne_28 & (~ IN2[24])  );
    wire logic pp_28_25;
    assign pp_28_25 = (select_e_28 & IN2[25] | select_2x_28 & IN2[24] | select_n2x_28 & (~ IN2[24]) | select_ne_28 & (~ IN2[25])  );
    wire logic pp_28_26;
    assign pp_28_26 = (select_e_28 & IN2[26] | select_2x_28 & IN2[25] | select_n2x_28 & (~ IN2[25]) | select_ne_28 & (~ IN2[26])  );
    wire logic pp_28_27;
    assign pp_28_27 = (select_e_28 & IN2[27] | select_2x_28 & IN2[26] | select_n2x_28 & (~ IN2[26]) | select_ne_28 & (~ IN2[27])  );
    wire logic pp_28_28;
    assign pp_28_28 = (select_e_28 & IN2[28] | select_2x_28 & IN2[27] | select_n2x_28 & (~ IN2[27]) | select_ne_28 & (~ IN2[28])  );
    wire logic pp_28_29;
    assign pp_28_29 = (select_e_28 & IN2[29] | select_2x_28 & IN2[28] | select_n2x_28 & (~ IN2[28]) | select_ne_28 & (~ IN2[29])  );
    wire logic pp_28_30;
    assign pp_28_30 = (select_e_28 & IN2[30] | select_2x_28 & IN2[29] | select_n2x_28 & (~ IN2[29]) | select_ne_28 & (~ IN2[30])  );
    wire logic pp_28_31;
    assign pp_28_31 = (select_e_28 & IN2[31] | select_2x_28 & IN2[30] | select_n2x_28 & (~ IN2[30]) | select_ne_28 & (~ IN2[31])  );
    wire logic pp_28_32;
    assign pp_28_32 = (select_e_28 & IN2[32] | select_2x_28 & IN2[31] | select_n2x_28 & (~ IN2[31]) | select_ne_28 & (~ IN2[32])  );
    wire logic pp_28_33;
    assign pp_28_33 = (select_e_28 & IN2[33] | select_2x_28 & IN2[32] | select_n2x_28 & (~ IN2[32]) | select_ne_28 & (~ IN2[33])  );
    wire logic pp_28_34;
    assign pp_28_34 = (select_e_28 & IN2[34] | select_2x_28 & IN2[33] | select_n2x_28 & (~ IN2[33]) | select_ne_28 & (~ IN2[34])  );
    wire logic pp_28_35;
    assign pp_28_35 = (select_e_28 & IN2[35] | select_2x_28 & IN2[34] | select_n2x_28 & (~ IN2[34]) | select_ne_28 & (~ IN2[35])  );
    wire logic pp_28_36;
    assign pp_28_36 = (select_e_28 & IN2[36] | select_2x_28 & IN2[35] | select_n2x_28 & (~ IN2[35]) | select_ne_28 & (~ IN2[36])  );
    wire logic pp_28_37;
    assign pp_28_37 = (select_e_28 & IN2[37] | select_2x_28 & IN2[36] | select_n2x_28 & (~ IN2[36]) | select_ne_28 & (~ IN2[37])  );
    wire logic pp_28_38;
    assign pp_28_38 = (select_e_28 & IN2[38] | select_2x_28 & IN2[37] | select_n2x_28 & (~ IN2[37]) | select_ne_28 & (~ IN2[38])  );
    wire logic pp_28_39;
    assign pp_28_39 = (select_e_28 & IN2[39] | select_2x_28 & IN2[38] | select_n2x_28 & (~ IN2[38]) | select_ne_28 & (~ IN2[39])  );
    wire logic pp_28_40;
    assign pp_28_40 = (select_e_28 & IN2[40] | select_2x_28 & IN2[39] | select_n2x_28 & (~ IN2[39]) | select_ne_28 & (~ IN2[40])  );
    wire logic pp_28_41;
    assign pp_28_41 = (select_e_28 & IN2[41] | select_2x_28 & IN2[40] | select_n2x_28 & (~ IN2[40]) | select_ne_28 & (~ IN2[41])  );
    wire logic pp_28_42;
    assign pp_28_42 = (select_e_28 & IN2[42] | select_2x_28 & IN2[41] | select_n2x_28 & (~ IN2[41]) | select_ne_28 & (~ IN2[42])  );
    wire logic pp_28_43;
    assign pp_28_43 = (select_e_28 & IN2[43] | select_2x_28 & IN2[42] | select_n2x_28 & (~ IN2[42]) | select_ne_28 & (~ IN2[43])  );
    wire logic pp_28_44;
    assign pp_28_44 = (select_e_28 & IN2[44] | select_2x_28 & IN2[43] | select_n2x_28 & (~ IN2[43]) | select_ne_28 & (~ IN2[44])  );
    wire logic pp_28_45;
    assign pp_28_45 = (select_e_28 & IN2[45] | select_2x_28 & IN2[44] | select_n2x_28 & (~ IN2[44]) | select_ne_28 & (~ IN2[45])  );
    wire logic pp_28_46;
    assign pp_28_46 = (select_e_28 & IN2[46] | select_2x_28 & IN2[45] | select_n2x_28 & (~ IN2[45]) | select_ne_28 & (~ IN2[46])  );
    wire logic pp_28_47;
    assign pp_28_47 = (select_e_28 & IN2[47] | select_2x_28 & IN2[46] | select_n2x_28 & (~ IN2[46]) | select_ne_28 & (~ IN2[47])  );
    wire logic pp_28_48;
    assign pp_28_48 = (select_e_28 & IN2[48] | select_2x_28 & IN2[47] | select_n2x_28 & (~ IN2[47]) | select_ne_28 & (~ IN2[48])  );
    wire logic pp_28_49;
    assign pp_28_49 = (select_e_28 & IN2[49] | select_2x_28 & IN2[48] | select_n2x_28 & (~ IN2[48]) | select_ne_28 & (~ IN2[49])  );
    wire logic pp_28_50;
    assign pp_28_50 = (select_e_28 & IN2[50] | select_2x_28 & IN2[49] | select_n2x_28 & (~ IN2[49]) | select_ne_28 & (~ IN2[50])  );
    wire logic pp_28_51;
    assign pp_28_51 = (select_e_28 & IN2[51] | select_2x_28 & IN2[50] | select_n2x_28 & (~ IN2[50]) | select_ne_28 & (~ IN2[51])  );
    wire logic pp_28_52;
    assign pp_28_52 = (select_e_28 & IN2[52] | select_2x_28 & IN2[51] | select_n2x_28 & (~ IN2[51]) | select_ne_28 & (~ IN2[52])  );
    wire logic pp_28_53;
    assign pp_28_53 = (select_e_28 & IN2[53] | select_2x_28 & IN2[52] | select_n2x_28 & (~ IN2[52]) | select_ne_28 & (~ IN2[53])  );
    wire logic pp_28_54;
    assign pp_28_54 = (select_e_28 & IN2[54] | select_2x_28 & IN2[53] | select_n2x_28 & (~ IN2[53]) | select_ne_28 & (~ IN2[54])  );
    wire logic pp_28_55;
    assign pp_28_55 = (select_e_28 & IN2[55] | select_2x_28 & IN2[54] | select_n2x_28 & (~ IN2[54]) | select_ne_28 & (~ IN2[55])  );
    wire logic pp_28_56;
    assign pp_28_56 = (select_e_28 & IN2[56] | select_2x_28 & IN2[55] | select_n2x_28 & (~ IN2[55]) | select_ne_28 & (~ IN2[56])  );
    wire logic pp_28_57;
    assign pp_28_57 = (select_e_28 & IN2[57] | select_2x_28 & IN2[56] | select_n2x_28 & (~ IN2[56]) | select_ne_28 & (~ IN2[57])  );
    wire logic pp_28_58;
    assign pp_28_58 = (select_e_28 & IN2[58] | select_2x_28 & IN2[57] | select_n2x_28 & (~ IN2[57]) | select_ne_28 & (~ IN2[58])  );
    wire logic pp_28_59;
    assign pp_28_59 = (select_e_28 & IN2[59] | select_2x_28 & IN2[58] | select_n2x_28 & (~ IN2[58]) | select_ne_28 & (~ IN2[59])  );
    wire logic pp_28_60;
    assign pp_28_60 = (select_e_28 & IN2[60] | select_2x_28 & IN2[59] | select_n2x_28 & (~ IN2[59]) | select_ne_28 & (~ IN2[60])  );
    wire logic pp_28_61;
    assign pp_28_61 = (select_e_28 & IN2[61] | select_2x_28 & IN2[60] | select_n2x_28 & (~ IN2[60]) | select_ne_28 & (~ IN2[61])  );
    wire logic pp_28_62;
    assign pp_28_62 = (select_e_28 & IN2[62] | select_2x_28 & IN2[61] | select_n2x_28 & (~ IN2[61]) | select_ne_28 & (~ IN2[62])  );
    wire logic pp_28_63;
    assign pp_28_63 = (select_e_28 & IN2[63] | select_2x_28 & IN2[62] | select_n2x_28 & (~ IN2[62]) | select_ne_28 & (~ IN2[63])  );
    wire logic pp_28_64;
    assign pp_28_64 = (select_e_28 & IN2[63] | select_2x_28 & IN2[63] | select_n2x_28 & (~ IN2[63]) | select_ne_28 & (~ IN2[63])  );
    wire logic pp_28_65;
    assign pp_28_65 = ~ (select_e_28 & IN2[63] | select_2x_28 & IN2[63] | select_n2x_28 & (~ IN2[63]) | select_ne_28 & (~ IN2[63])  );
    assign tcomp28 = select_ne_28 | select_n2x_28;
    
    // Signed Booth Radix-4 Partial Products Row 30
    wire logic select_e_29, select_ne_29, select_2x_29, tcomp29, select_n2x_29;
    assign select_e_29 = ((~ IN1[59]) & (IN1[58] ^ IN1[57]));
    assign select_ne_29 = IN1[59] &  (IN1[58] ^ IN1[57]);
    assign select_2x_29 = (~ IN1[59]) & IN1[58] & IN1[57];
    assign select_n2x_29 = IN1[59] & (~ IN1[58]) & (~ IN1[57]);
    wire logic pp_29_0;
    assign pp_29_0 = (select_e_29 & IN2[0] | select_2x_29 & 1'b0 | select_n2x_29 & 1'b1 | select_ne_29 & (~ IN2[0])  );
    wire logic pp_29_1;
    assign pp_29_1 = (select_e_29 & IN2[1] | select_2x_29 & IN2[0] | select_n2x_29 & (~ IN2[0]) | select_ne_29 & (~ IN2[1])  );
    wire logic pp_29_2;
    assign pp_29_2 = (select_e_29 & IN2[2] | select_2x_29 & IN2[1] | select_n2x_29 & (~ IN2[1]) | select_ne_29 & (~ IN2[2])  );
    wire logic pp_29_3;
    assign pp_29_3 = (select_e_29 & IN2[3] | select_2x_29 & IN2[2] | select_n2x_29 & (~ IN2[2]) | select_ne_29 & (~ IN2[3])  );
    wire logic pp_29_4;
    assign pp_29_4 = (select_e_29 & IN2[4] | select_2x_29 & IN2[3] | select_n2x_29 & (~ IN2[3]) | select_ne_29 & (~ IN2[4])  );
    wire logic pp_29_5;
    assign pp_29_5 = (select_e_29 & IN2[5] | select_2x_29 & IN2[4] | select_n2x_29 & (~ IN2[4]) | select_ne_29 & (~ IN2[5])  );
    wire logic pp_29_6;
    assign pp_29_6 = (select_e_29 & IN2[6] | select_2x_29 & IN2[5] | select_n2x_29 & (~ IN2[5]) | select_ne_29 & (~ IN2[6])  );
    wire logic pp_29_7;
    assign pp_29_7 = (select_e_29 & IN2[7] | select_2x_29 & IN2[6] | select_n2x_29 & (~ IN2[6]) | select_ne_29 & (~ IN2[7])  );
    wire logic pp_29_8;
    assign pp_29_8 = (select_e_29 & IN2[8] | select_2x_29 & IN2[7] | select_n2x_29 & (~ IN2[7]) | select_ne_29 & (~ IN2[8])  );
    wire logic pp_29_9;
    assign pp_29_9 = (select_e_29 & IN2[9] | select_2x_29 & IN2[8] | select_n2x_29 & (~ IN2[8]) | select_ne_29 & (~ IN2[9])  );
    wire logic pp_29_10;
    assign pp_29_10 = (select_e_29 & IN2[10] | select_2x_29 & IN2[9] | select_n2x_29 & (~ IN2[9]) | select_ne_29 & (~ IN2[10])  );
    wire logic pp_29_11;
    assign pp_29_11 = (select_e_29 & IN2[11] | select_2x_29 & IN2[10] | select_n2x_29 & (~ IN2[10]) | select_ne_29 & (~ IN2[11])  );
    wire logic pp_29_12;
    assign pp_29_12 = (select_e_29 & IN2[12] | select_2x_29 & IN2[11] | select_n2x_29 & (~ IN2[11]) | select_ne_29 & (~ IN2[12])  );
    wire logic pp_29_13;
    assign pp_29_13 = (select_e_29 & IN2[13] | select_2x_29 & IN2[12] | select_n2x_29 & (~ IN2[12]) | select_ne_29 & (~ IN2[13])  );
    wire logic pp_29_14;
    assign pp_29_14 = (select_e_29 & IN2[14] | select_2x_29 & IN2[13] | select_n2x_29 & (~ IN2[13]) | select_ne_29 & (~ IN2[14])  );
    wire logic pp_29_15;
    assign pp_29_15 = (select_e_29 & IN2[15] | select_2x_29 & IN2[14] | select_n2x_29 & (~ IN2[14]) | select_ne_29 & (~ IN2[15])  );
    wire logic pp_29_16;
    assign pp_29_16 = (select_e_29 & IN2[16] | select_2x_29 & IN2[15] | select_n2x_29 & (~ IN2[15]) | select_ne_29 & (~ IN2[16])  );
    wire logic pp_29_17;
    assign pp_29_17 = (select_e_29 & IN2[17] | select_2x_29 & IN2[16] | select_n2x_29 & (~ IN2[16]) | select_ne_29 & (~ IN2[17])  );
    wire logic pp_29_18;
    assign pp_29_18 = (select_e_29 & IN2[18] | select_2x_29 & IN2[17] | select_n2x_29 & (~ IN2[17]) | select_ne_29 & (~ IN2[18])  );
    wire logic pp_29_19;
    assign pp_29_19 = (select_e_29 & IN2[19] | select_2x_29 & IN2[18] | select_n2x_29 & (~ IN2[18]) | select_ne_29 & (~ IN2[19])  );
    wire logic pp_29_20;
    assign pp_29_20 = (select_e_29 & IN2[20] | select_2x_29 & IN2[19] | select_n2x_29 & (~ IN2[19]) | select_ne_29 & (~ IN2[20])  );
    wire logic pp_29_21;
    assign pp_29_21 = (select_e_29 & IN2[21] | select_2x_29 & IN2[20] | select_n2x_29 & (~ IN2[20]) | select_ne_29 & (~ IN2[21])  );
    wire logic pp_29_22;
    assign pp_29_22 = (select_e_29 & IN2[22] | select_2x_29 & IN2[21] | select_n2x_29 & (~ IN2[21]) | select_ne_29 & (~ IN2[22])  );
    wire logic pp_29_23;
    assign pp_29_23 = (select_e_29 & IN2[23] | select_2x_29 & IN2[22] | select_n2x_29 & (~ IN2[22]) | select_ne_29 & (~ IN2[23])  );
    wire logic pp_29_24;
    assign pp_29_24 = (select_e_29 & IN2[24] | select_2x_29 & IN2[23] | select_n2x_29 & (~ IN2[23]) | select_ne_29 & (~ IN2[24])  );
    wire logic pp_29_25;
    assign pp_29_25 = (select_e_29 & IN2[25] | select_2x_29 & IN2[24] | select_n2x_29 & (~ IN2[24]) | select_ne_29 & (~ IN2[25])  );
    wire logic pp_29_26;
    assign pp_29_26 = (select_e_29 & IN2[26] | select_2x_29 & IN2[25] | select_n2x_29 & (~ IN2[25]) | select_ne_29 & (~ IN2[26])  );
    wire logic pp_29_27;
    assign pp_29_27 = (select_e_29 & IN2[27] | select_2x_29 & IN2[26] | select_n2x_29 & (~ IN2[26]) | select_ne_29 & (~ IN2[27])  );
    wire logic pp_29_28;
    assign pp_29_28 = (select_e_29 & IN2[28] | select_2x_29 & IN2[27] | select_n2x_29 & (~ IN2[27]) | select_ne_29 & (~ IN2[28])  );
    wire logic pp_29_29;
    assign pp_29_29 = (select_e_29 & IN2[29] | select_2x_29 & IN2[28] | select_n2x_29 & (~ IN2[28]) | select_ne_29 & (~ IN2[29])  );
    wire logic pp_29_30;
    assign pp_29_30 = (select_e_29 & IN2[30] | select_2x_29 & IN2[29] | select_n2x_29 & (~ IN2[29]) | select_ne_29 & (~ IN2[30])  );
    wire logic pp_29_31;
    assign pp_29_31 = (select_e_29 & IN2[31] | select_2x_29 & IN2[30] | select_n2x_29 & (~ IN2[30]) | select_ne_29 & (~ IN2[31])  );
    wire logic pp_29_32;
    assign pp_29_32 = (select_e_29 & IN2[32] | select_2x_29 & IN2[31] | select_n2x_29 & (~ IN2[31]) | select_ne_29 & (~ IN2[32])  );
    wire logic pp_29_33;
    assign pp_29_33 = (select_e_29 & IN2[33] | select_2x_29 & IN2[32] | select_n2x_29 & (~ IN2[32]) | select_ne_29 & (~ IN2[33])  );
    wire logic pp_29_34;
    assign pp_29_34 = (select_e_29 & IN2[34] | select_2x_29 & IN2[33] | select_n2x_29 & (~ IN2[33]) | select_ne_29 & (~ IN2[34])  );
    wire logic pp_29_35;
    assign pp_29_35 = (select_e_29 & IN2[35] | select_2x_29 & IN2[34] | select_n2x_29 & (~ IN2[34]) | select_ne_29 & (~ IN2[35])  );
    wire logic pp_29_36;
    assign pp_29_36 = (select_e_29 & IN2[36] | select_2x_29 & IN2[35] | select_n2x_29 & (~ IN2[35]) | select_ne_29 & (~ IN2[36])  );
    wire logic pp_29_37;
    assign pp_29_37 = (select_e_29 & IN2[37] | select_2x_29 & IN2[36] | select_n2x_29 & (~ IN2[36]) | select_ne_29 & (~ IN2[37])  );
    wire logic pp_29_38;
    assign pp_29_38 = (select_e_29 & IN2[38] | select_2x_29 & IN2[37] | select_n2x_29 & (~ IN2[37]) | select_ne_29 & (~ IN2[38])  );
    wire logic pp_29_39;
    assign pp_29_39 = (select_e_29 & IN2[39] | select_2x_29 & IN2[38] | select_n2x_29 & (~ IN2[38]) | select_ne_29 & (~ IN2[39])  );
    wire logic pp_29_40;
    assign pp_29_40 = (select_e_29 & IN2[40] | select_2x_29 & IN2[39] | select_n2x_29 & (~ IN2[39]) | select_ne_29 & (~ IN2[40])  );
    wire logic pp_29_41;
    assign pp_29_41 = (select_e_29 & IN2[41] | select_2x_29 & IN2[40] | select_n2x_29 & (~ IN2[40]) | select_ne_29 & (~ IN2[41])  );
    wire logic pp_29_42;
    assign pp_29_42 = (select_e_29 & IN2[42] | select_2x_29 & IN2[41] | select_n2x_29 & (~ IN2[41]) | select_ne_29 & (~ IN2[42])  );
    wire logic pp_29_43;
    assign pp_29_43 = (select_e_29 & IN2[43] | select_2x_29 & IN2[42] | select_n2x_29 & (~ IN2[42]) | select_ne_29 & (~ IN2[43])  );
    wire logic pp_29_44;
    assign pp_29_44 = (select_e_29 & IN2[44] | select_2x_29 & IN2[43] | select_n2x_29 & (~ IN2[43]) | select_ne_29 & (~ IN2[44])  );
    wire logic pp_29_45;
    assign pp_29_45 = (select_e_29 & IN2[45] | select_2x_29 & IN2[44] | select_n2x_29 & (~ IN2[44]) | select_ne_29 & (~ IN2[45])  );
    wire logic pp_29_46;
    assign pp_29_46 = (select_e_29 & IN2[46] | select_2x_29 & IN2[45] | select_n2x_29 & (~ IN2[45]) | select_ne_29 & (~ IN2[46])  );
    wire logic pp_29_47;
    assign pp_29_47 = (select_e_29 & IN2[47] | select_2x_29 & IN2[46] | select_n2x_29 & (~ IN2[46]) | select_ne_29 & (~ IN2[47])  );
    wire logic pp_29_48;
    assign pp_29_48 = (select_e_29 & IN2[48] | select_2x_29 & IN2[47] | select_n2x_29 & (~ IN2[47]) | select_ne_29 & (~ IN2[48])  );
    wire logic pp_29_49;
    assign pp_29_49 = (select_e_29 & IN2[49] | select_2x_29 & IN2[48] | select_n2x_29 & (~ IN2[48]) | select_ne_29 & (~ IN2[49])  );
    wire logic pp_29_50;
    assign pp_29_50 = (select_e_29 & IN2[50] | select_2x_29 & IN2[49] | select_n2x_29 & (~ IN2[49]) | select_ne_29 & (~ IN2[50])  );
    wire logic pp_29_51;
    assign pp_29_51 = (select_e_29 & IN2[51] | select_2x_29 & IN2[50] | select_n2x_29 & (~ IN2[50]) | select_ne_29 & (~ IN2[51])  );
    wire logic pp_29_52;
    assign pp_29_52 = (select_e_29 & IN2[52] | select_2x_29 & IN2[51] | select_n2x_29 & (~ IN2[51]) | select_ne_29 & (~ IN2[52])  );
    wire logic pp_29_53;
    assign pp_29_53 = (select_e_29 & IN2[53] | select_2x_29 & IN2[52] | select_n2x_29 & (~ IN2[52]) | select_ne_29 & (~ IN2[53])  );
    wire logic pp_29_54;
    assign pp_29_54 = (select_e_29 & IN2[54] | select_2x_29 & IN2[53] | select_n2x_29 & (~ IN2[53]) | select_ne_29 & (~ IN2[54])  );
    wire logic pp_29_55;
    assign pp_29_55 = (select_e_29 & IN2[55] | select_2x_29 & IN2[54] | select_n2x_29 & (~ IN2[54]) | select_ne_29 & (~ IN2[55])  );
    wire logic pp_29_56;
    assign pp_29_56 = (select_e_29 & IN2[56] | select_2x_29 & IN2[55] | select_n2x_29 & (~ IN2[55]) | select_ne_29 & (~ IN2[56])  );
    wire logic pp_29_57;
    assign pp_29_57 = (select_e_29 & IN2[57] | select_2x_29 & IN2[56] | select_n2x_29 & (~ IN2[56]) | select_ne_29 & (~ IN2[57])  );
    wire logic pp_29_58;
    assign pp_29_58 = (select_e_29 & IN2[58] | select_2x_29 & IN2[57] | select_n2x_29 & (~ IN2[57]) | select_ne_29 & (~ IN2[58])  );
    wire logic pp_29_59;
    assign pp_29_59 = (select_e_29 & IN2[59] | select_2x_29 & IN2[58] | select_n2x_29 & (~ IN2[58]) | select_ne_29 & (~ IN2[59])  );
    wire logic pp_29_60;
    assign pp_29_60 = (select_e_29 & IN2[60] | select_2x_29 & IN2[59] | select_n2x_29 & (~ IN2[59]) | select_ne_29 & (~ IN2[60])  );
    wire logic pp_29_61;
    assign pp_29_61 = (select_e_29 & IN2[61] | select_2x_29 & IN2[60] | select_n2x_29 & (~ IN2[60]) | select_ne_29 & (~ IN2[61])  );
    wire logic pp_29_62;
    assign pp_29_62 = (select_e_29 & IN2[62] | select_2x_29 & IN2[61] | select_n2x_29 & (~ IN2[61]) | select_ne_29 & (~ IN2[62])  );
    wire logic pp_29_63;
    assign pp_29_63 = (select_e_29 & IN2[63] | select_2x_29 & IN2[62] | select_n2x_29 & (~ IN2[62]) | select_ne_29 & (~ IN2[63])  );
    wire logic pp_29_64;
    assign pp_29_64 = (select_e_29 & IN2[63] | select_2x_29 & IN2[63] | select_n2x_29 & (~ IN2[63]) | select_ne_29 & (~ IN2[63])  );
    wire logic pp_29_65;
    assign pp_29_65 = ~ (select_e_29 & IN2[63] | select_2x_29 & IN2[63] | select_n2x_29 & (~ IN2[63]) | select_ne_29 & (~ IN2[63])  );
    assign tcomp29 = select_ne_29 | select_n2x_29;
    
    // Signed Booth Radix-4 Partial Products Row 31
    wire logic select_e_30, select_ne_30, select_2x_30, tcomp30, select_n2x_30;
    assign select_e_30 = ((~ IN1[61]) & (IN1[60] ^ IN1[59]));
    assign select_ne_30 = IN1[61] &  (IN1[60] ^ IN1[59]);
    assign select_2x_30 = (~ IN1[61]) & IN1[60] & IN1[59];
    assign select_n2x_30 = IN1[61] & (~ IN1[60]) & (~ IN1[59]);
    wire logic pp_30_0;
    assign pp_30_0 = (select_e_30 & IN2[0] | select_2x_30 & 1'b0 | select_n2x_30 & 1'b1 | select_ne_30 & (~ IN2[0])  );
    wire logic pp_30_1;
    assign pp_30_1 = (select_e_30 & IN2[1] | select_2x_30 & IN2[0] | select_n2x_30 & (~ IN2[0]) | select_ne_30 & (~ IN2[1])  );
    wire logic pp_30_2;
    assign pp_30_2 = (select_e_30 & IN2[2] | select_2x_30 & IN2[1] | select_n2x_30 & (~ IN2[1]) | select_ne_30 & (~ IN2[2])  );
    wire logic pp_30_3;
    assign pp_30_3 = (select_e_30 & IN2[3] | select_2x_30 & IN2[2] | select_n2x_30 & (~ IN2[2]) | select_ne_30 & (~ IN2[3])  );
    wire logic pp_30_4;
    assign pp_30_4 = (select_e_30 & IN2[4] | select_2x_30 & IN2[3] | select_n2x_30 & (~ IN2[3]) | select_ne_30 & (~ IN2[4])  );
    wire logic pp_30_5;
    assign pp_30_5 = (select_e_30 & IN2[5] | select_2x_30 & IN2[4] | select_n2x_30 & (~ IN2[4]) | select_ne_30 & (~ IN2[5])  );
    wire logic pp_30_6;
    assign pp_30_6 = (select_e_30 & IN2[6] | select_2x_30 & IN2[5] | select_n2x_30 & (~ IN2[5]) | select_ne_30 & (~ IN2[6])  );
    wire logic pp_30_7;
    assign pp_30_7 = (select_e_30 & IN2[7] | select_2x_30 & IN2[6] | select_n2x_30 & (~ IN2[6]) | select_ne_30 & (~ IN2[7])  );
    wire logic pp_30_8;
    assign pp_30_8 = (select_e_30 & IN2[8] | select_2x_30 & IN2[7] | select_n2x_30 & (~ IN2[7]) | select_ne_30 & (~ IN2[8])  );
    wire logic pp_30_9;
    assign pp_30_9 = (select_e_30 & IN2[9] | select_2x_30 & IN2[8] | select_n2x_30 & (~ IN2[8]) | select_ne_30 & (~ IN2[9])  );
    wire logic pp_30_10;
    assign pp_30_10 = (select_e_30 & IN2[10] | select_2x_30 & IN2[9] | select_n2x_30 & (~ IN2[9]) | select_ne_30 & (~ IN2[10])  );
    wire logic pp_30_11;
    assign pp_30_11 = (select_e_30 & IN2[11] | select_2x_30 & IN2[10] | select_n2x_30 & (~ IN2[10]) | select_ne_30 & (~ IN2[11])  );
    wire logic pp_30_12;
    assign pp_30_12 = (select_e_30 & IN2[12] | select_2x_30 & IN2[11] | select_n2x_30 & (~ IN2[11]) | select_ne_30 & (~ IN2[12])  );
    wire logic pp_30_13;
    assign pp_30_13 = (select_e_30 & IN2[13] | select_2x_30 & IN2[12] | select_n2x_30 & (~ IN2[12]) | select_ne_30 & (~ IN2[13])  );
    wire logic pp_30_14;
    assign pp_30_14 = (select_e_30 & IN2[14] | select_2x_30 & IN2[13] | select_n2x_30 & (~ IN2[13]) | select_ne_30 & (~ IN2[14])  );
    wire logic pp_30_15;
    assign pp_30_15 = (select_e_30 & IN2[15] | select_2x_30 & IN2[14] | select_n2x_30 & (~ IN2[14]) | select_ne_30 & (~ IN2[15])  );
    wire logic pp_30_16;
    assign pp_30_16 = (select_e_30 & IN2[16] | select_2x_30 & IN2[15] | select_n2x_30 & (~ IN2[15]) | select_ne_30 & (~ IN2[16])  );
    wire logic pp_30_17;
    assign pp_30_17 = (select_e_30 & IN2[17] | select_2x_30 & IN2[16] | select_n2x_30 & (~ IN2[16]) | select_ne_30 & (~ IN2[17])  );
    wire logic pp_30_18;
    assign pp_30_18 = (select_e_30 & IN2[18] | select_2x_30 & IN2[17] | select_n2x_30 & (~ IN2[17]) | select_ne_30 & (~ IN2[18])  );
    wire logic pp_30_19;
    assign pp_30_19 = (select_e_30 & IN2[19] | select_2x_30 & IN2[18] | select_n2x_30 & (~ IN2[18]) | select_ne_30 & (~ IN2[19])  );
    wire logic pp_30_20;
    assign pp_30_20 = (select_e_30 & IN2[20] | select_2x_30 & IN2[19] | select_n2x_30 & (~ IN2[19]) | select_ne_30 & (~ IN2[20])  );
    wire logic pp_30_21;
    assign pp_30_21 = (select_e_30 & IN2[21] | select_2x_30 & IN2[20] | select_n2x_30 & (~ IN2[20]) | select_ne_30 & (~ IN2[21])  );
    wire logic pp_30_22;
    assign pp_30_22 = (select_e_30 & IN2[22] | select_2x_30 & IN2[21] | select_n2x_30 & (~ IN2[21]) | select_ne_30 & (~ IN2[22])  );
    wire logic pp_30_23;
    assign pp_30_23 = (select_e_30 & IN2[23] | select_2x_30 & IN2[22] | select_n2x_30 & (~ IN2[22]) | select_ne_30 & (~ IN2[23])  );
    wire logic pp_30_24;
    assign pp_30_24 = (select_e_30 & IN2[24] | select_2x_30 & IN2[23] | select_n2x_30 & (~ IN2[23]) | select_ne_30 & (~ IN2[24])  );
    wire logic pp_30_25;
    assign pp_30_25 = (select_e_30 & IN2[25] | select_2x_30 & IN2[24] | select_n2x_30 & (~ IN2[24]) | select_ne_30 & (~ IN2[25])  );
    wire logic pp_30_26;
    assign pp_30_26 = (select_e_30 & IN2[26] | select_2x_30 & IN2[25] | select_n2x_30 & (~ IN2[25]) | select_ne_30 & (~ IN2[26])  );
    wire logic pp_30_27;
    assign pp_30_27 = (select_e_30 & IN2[27] | select_2x_30 & IN2[26] | select_n2x_30 & (~ IN2[26]) | select_ne_30 & (~ IN2[27])  );
    wire logic pp_30_28;
    assign pp_30_28 = (select_e_30 & IN2[28] | select_2x_30 & IN2[27] | select_n2x_30 & (~ IN2[27]) | select_ne_30 & (~ IN2[28])  );
    wire logic pp_30_29;
    assign pp_30_29 = (select_e_30 & IN2[29] | select_2x_30 & IN2[28] | select_n2x_30 & (~ IN2[28]) | select_ne_30 & (~ IN2[29])  );
    wire logic pp_30_30;
    assign pp_30_30 = (select_e_30 & IN2[30] | select_2x_30 & IN2[29] | select_n2x_30 & (~ IN2[29]) | select_ne_30 & (~ IN2[30])  );
    wire logic pp_30_31;
    assign pp_30_31 = (select_e_30 & IN2[31] | select_2x_30 & IN2[30] | select_n2x_30 & (~ IN2[30]) | select_ne_30 & (~ IN2[31])  );
    wire logic pp_30_32;
    assign pp_30_32 = (select_e_30 & IN2[32] | select_2x_30 & IN2[31] | select_n2x_30 & (~ IN2[31]) | select_ne_30 & (~ IN2[32])  );
    wire logic pp_30_33;
    assign pp_30_33 = (select_e_30 & IN2[33] | select_2x_30 & IN2[32] | select_n2x_30 & (~ IN2[32]) | select_ne_30 & (~ IN2[33])  );
    wire logic pp_30_34;
    assign pp_30_34 = (select_e_30 & IN2[34] | select_2x_30 & IN2[33] | select_n2x_30 & (~ IN2[33]) | select_ne_30 & (~ IN2[34])  );
    wire logic pp_30_35;
    assign pp_30_35 = (select_e_30 & IN2[35] | select_2x_30 & IN2[34] | select_n2x_30 & (~ IN2[34]) | select_ne_30 & (~ IN2[35])  );
    wire logic pp_30_36;
    assign pp_30_36 = (select_e_30 & IN2[36] | select_2x_30 & IN2[35] | select_n2x_30 & (~ IN2[35]) | select_ne_30 & (~ IN2[36])  );
    wire logic pp_30_37;
    assign pp_30_37 = (select_e_30 & IN2[37] | select_2x_30 & IN2[36] | select_n2x_30 & (~ IN2[36]) | select_ne_30 & (~ IN2[37])  );
    wire logic pp_30_38;
    assign pp_30_38 = (select_e_30 & IN2[38] | select_2x_30 & IN2[37] | select_n2x_30 & (~ IN2[37]) | select_ne_30 & (~ IN2[38])  );
    wire logic pp_30_39;
    assign pp_30_39 = (select_e_30 & IN2[39] | select_2x_30 & IN2[38] | select_n2x_30 & (~ IN2[38]) | select_ne_30 & (~ IN2[39])  );
    wire logic pp_30_40;
    assign pp_30_40 = (select_e_30 & IN2[40] | select_2x_30 & IN2[39] | select_n2x_30 & (~ IN2[39]) | select_ne_30 & (~ IN2[40])  );
    wire logic pp_30_41;
    assign pp_30_41 = (select_e_30 & IN2[41] | select_2x_30 & IN2[40] | select_n2x_30 & (~ IN2[40]) | select_ne_30 & (~ IN2[41])  );
    wire logic pp_30_42;
    assign pp_30_42 = (select_e_30 & IN2[42] | select_2x_30 & IN2[41] | select_n2x_30 & (~ IN2[41]) | select_ne_30 & (~ IN2[42])  );
    wire logic pp_30_43;
    assign pp_30_43 = (select_e_30 & IN2[43] | select_2x_30 & IN2[42] | select_n2x_30 & (~ IN2[42]) | select_ne_30 & (~ IN2[43])  );
    wire logic pp_30_44;
    assign pp_30_44 = (select_e_30 & IN2[44] | select_2x_30 & IN2[43] | select_n2x_30 & (~ IN2[43]) | select_ne_30 & (~ IN2[44])  );
    wire logic pp_30_45;
    assign pp_30_45 = (select_e_30 & IN2[45] | select_2x_30 & IN2[44] | select_n2x_30 & (~ IN2[44]) | select_ne_30 & (~ IN2[45])  );
    wire logic pp_30_46;
    assign pp_30_46 = (select_e_30 & IN2[46] | select_2x_30 & IN2[45] | select_n2x_30 & (~ IN2[45]) | select_ne_30 & (~ IN2[46])  );
    wire logic pp_30_47;
    assign pp_30_47 = (select_e_30 & IN2[47] | select_2x_30 & IN2[46] | select_n2x_30 & (~ IN2[46]) | select_ne_30 & (~ IN2[47])  );
    wire logic pp_30_48;
    assign pp_30_48 = (select_e_30 & IN2[48] | select_2x_30 & IN2[47] | select_n2x_30 & (~ IN2[47]) | select_ne_30 & (~ IN2[48])  );
    wire logic pp_30_49;
    assign pp_30_49 = (select_e_30 & IN2[49] | select_2x_30 & IN2[48] | select_n2x_30 & (~ IN2[48]) | select_ne_30 & (~ IN2[49])  );
    wire logic pp_30_50;
    assign pp_30_50 = (select_e_30 & IN2[50] | select_2x_30 & IN2[49] | select_n2x_30 & (~ IN2[49]) | select_ne_30 & (~ IN2[50])  );
    wire logic pp_30_51;
    assign pp_30_51 = (select_e_30 & IN2[51] | select_2x_30 & IN2[50] | select_n2x_30 & (~ IN2[50]) | select_ne_30 & (~ IN2[51])  );
    wire logic pp_30_52;
    assign pp_30_52 = (select_e_30 & IN2[52] | select_2x_30 & IN2[51] | select_n2x_30 & (~ IN2[51]) | select_ne_30 & (~ IN2[52])  );
    wire logic pp_30_53;
    assign pp_30_53 = (select_e_30 & IN2[53] | select_2x_30 & IN2[52] | select_n2x_30 & (~ IN2[52]) | select_ne_30 & (~ IN2[53])  );
    wire logic pp_30_54;
    assign pp_30_54 = (select_e_30 & IN2[54] | select_2x_30 & IN2[53] | select_n2x_30 & (~ IN2[53]) | select_ne_30 & (~ IN2[54])  );
    wire logic pp_30_55;
    assign pp_30_55 = (select_e_30 & IN2[55] | select_2x_30 & IN2[54] | select_n2x_30 & (~ IN2[54]) | select_ne_30 & (~ IN2[55])  );
    wire logic pp_30_56;
    assign pp_30_56 = (select_e_30 & IN2[56] | select_2x_30 & IN2[55] | select_n2x_30 & (~ IN2[55]) | select_ne_30 & (~ IN2[56])  );
    wire logic pp_30_57;
    assign pp_30_57 = (select_e_30 & IN2[57] | select_2x_30 & IN2[56] | select_n2x_30 & (~ IN2[56]) | select_ne_30 & (~ IN2[57])  );
    wire logic pp_30_58;
    assign pp_30_58 = (select_e_30 & IN2[58] | select_2x_30 & IN2[57] | select_n2x_30 & (~ IN2[57]) | select_ne_30 & (~ IN2[58])  );
    wire logic pp_30_59;
    assign pp_30_59 = (select_e_30 & IN2[59] | select_2x_30 & IN2[58] | select_n2x_30 & (~ IN2[58]) | select_ne_30 & (~ IN2[59])  );
    wire logic pp_30_60;
    assign pp_30_60 = (select_e_30 & IN2[60] | select_2x_30 & IN2[59] | select_n2x_30 & (~ IN2[59]) | select_ne_30 & (~ IN2[60])  );
    wire logic pp_30_61;
    assign pp_30_61 = (select_e_30 & IN2[61] | select_2x_30 & IN2[60] | select_n2x_30 & (~ IN2[60]) | select_ne_30 & (~ IN2[61])  );
    wire logic pp_30_62;
    assign pp_30_62 = (select_e_30 & IN2[62] | select_2x_30 & IN2[61] | select_n2x_30 & (~ IN2[61]) | select_ne_30 & (~ IN2[62])  );
    wire logic pp_30_63;
    assign pp_30_63 = (select_e_30 & IN2[63] | select_2x_30 & IN2[62] | select_n2x_30 & (~ IN2[62]) | select_ne_30 & (~ IN2[63])  );
    wire logic pp_30_64;
    assign pp_30_64 = (select_e_30 & IN2[63] | select_2x_30 & IN2[63] | select_n2x_30 & (~ IN2[63]) | select_ne_30 & (~ IN2[63])  );
    wire logic pp_30_65;
    assign pp_30_65 = ~ (select_e_30 & IN2[63] | select_2x_30 & IN2[63] | select_n2x_30 & (~ IN2[63]) | select_ne_30 & (~ IN2[63])  );
    assign tcomp30 = select_ne_30 | select_n2x_30;
    
    // Signed Booth Radix-4 Partial Products Row 32
    wire logic select_e_31, select_ne_31, select_2x_31, tcomp31, select_n2x_31;
    assign select_e_31 = ((~ IN1[63]) & (IN1[62] ^ IN1[61]));
    assign select_ne_31 = IN1[63] &  (IN1[62] ^ IN1[61]);
    assign select_2x_31 = (~ IN1[63]) & IN1[62] & IN1[61];
    assign select_n2x_31 = IN1[63] & (~ IN1[62]) & (~ IN1[61]);
    wire logic pp_31_0;
    assign pp_31_0 = (select_e_31 & IN2[0] | select_2x_31 & 1'b0 | select_n2x_31 & 1'b1 | select_ne_31 & (~ IN2[0])  );
    wire logic pp_31_1;
    assign pp_31_1 = (select_e_31 & IN2[1] | select_2x_31 & IN2[0] | select_n2x_31 & (~ IN2[0]) | select_ne_31 & (~ IN2[1])  );
    wire logic pp_31_2;
    assign pp_31_2 = (select_e_31 & IN2[2] | select_2x_31 & IN2[1] | select_n2x_31 & (~ IN2[1]) | select_ne_31 & (~ IN2[2])  );
    wire logic pp_31_3;
    assign pp_31_3 = (select_e_31 & IN2[3] | select_2x_31 & IN2[2] | select_n2x_31 & (~ IN2[2]) | select_ne_31 & (~ IN2[3])  );
    wire logic pp_31_4;
    assign pp_31_4 = (select_e_31 & IN2[4] | select_2x_31 & IN2[3] | select_n2x_31 & (~ IN2[3]) | select_ne_31 & (~ IN2[4])  );
    wire logic pp_31_5;
    assign pp_31_5 = (select_e_31 & IN2[5] | select_2x_31 & IN2[4] | select_n2x_31 & (~ IN2[4]) | select_ne_31 & (~ IN2[5])  );
    wire logic pp_31_6;
    assign pp_31_6 = (select_e_31 & IN2[6] | select_2x_31 & IN2[5] | select_n2x_31 & (~ IN2[5]) | select_ne_31 & (~ IN2[6])  );
    wire logic pp_31_7;
    assign pp_31_7 = (select_e_31 & IN2[7] | select_2x_31 & IN2[6] | select_n2x_31 & (~ IN2[6]) | select_ne_31 & (~ IN2[7])  );
    wire logic pp_31_8;
    assign pp_31_8 = (select_e_31 & IN2[8] | select_2x_31 & IN2[7] | select_n2x_31 & (~ IN2[7]) | select_ne_31 & (~ IN2[8])  );
    wire logic pp_31_9;
    assign pp_31_9 = (select_e_31 & IN2[9] | select_2x_31 & IN2[8] | select_n2x_31 & (~ IN2[8]) | select_ne_31 & (~ IN2[9])  );
    wire logic pp_31_10;
    assign pp_31_10 = (select_e_31 & IN2[10] | select_2x_31 & IN2[9] | select_n2x_31 & (~ IN2[9]) | select_ne_31 & (~ IN2[10])  );
    wire logic pp_31_11;
    assign pp_31_11 = (select_e_31 & IN2[11] | select_2x_31 & IN2[10] | select_n2x_31 & (~ IN2[10]) | select_ne_31 & (~ IN2[11])  );
    wire logic pp_31_12;
    assign pp_31_12 = (select_e_31 & IN2[12] | select_2x_31 & IN2[11] | select_n2x_31 & (~ IN2[11]) | select_ne_31 & (~ IN2[12])  );
    wire logic pp_31_13;
    assign pp_31_13 = (select_e_31 & IN2[13] | select_2x_31 & IN2[12] | select_n2x_31 & (~ IN2[12]) | select_ne_31 & (~ IN2[13])  );
    wire logic pp_31_14;
    assign pp_31_14 = (select_e_31 & IN2[14] | select_2x_31 & IN2[13] | select_n2x_31 & (~ IN2[13]) | select_ne_31 & (~ IN2[14])  );
    wire logic pp_31_15;
    assign pp_31_15 = (select_e_31 & IN2[15] | select_2x_31 & IN2[14] | select_n2x_31 & (~ IN2[14]) | select_ne_31 & (~ IN2[15])  );
    wire logic pp_31_16;
    assign pp_31_16 = (select_e_31 & IN2[16] | select_2x_31 & IN2[15] | select_n2x_31 & (~ IN2[15]) | select_ne_31 & (~ IN2[16])  );
    wire logic pp_31_17;
    assign pp_31_17 = (select_e_31 & IN2[17] | select_2x_31 & IN2[16] | select_n2x_31 & (~ IN2[16]) | select_ne_31 & (~ IN2[17])  );
    wire logic pp_31_18;
    assign pp_31_18 = (select_e_31 & IN2[18] | select_2x_31 & IN2[17] | select_n2x_31 & (~ IN2[17]) | select_ne_31 & (~ IN2[18])  );
    wire logic pp_31_19;
    assign pp_31_19 = (select_e_31 & IN2[19] | select_2x_31 & IN2[18] | select_n2x_31 & (~ IN2[18]) | select_ne_31 & (~ IN2[19])  );
    wire logic pp_31_20;
    assign pp_31_20 = (select_e_31 & IN2[20] | select_2x_31 & IN2[19] | select_n2x_31 & (~ IN2[19]) | select_ne_31 & (~ IN2[20])  );
    wire logic pp_31_21;
    assign pp_31_21 = (select_e_31 & IN2[21] | select_2x_31 & IN2[20] | select_n2x_31 & (~ IN2[20]) | select_ne_31 & (~ IN2[21])  );
    wire logic pp_31_22;
    assign pp_31_22 = (select_e_31 & IN2[22] | select_2x_31 & IN2[21] | select_n2x_31 & (~ IN2[21]) | select_ne_31 & (~ IN2[22])  );
    wire logic pp_31_23;
    assign pp_31_23 = (select_e_31 & IN2[23] | select_2x_31 & IN2[22] | select_n2x_31 & (~ IN2[22]) | select_ne_31 & (~ IN2[23])  );
    wire logic pp_31_24;
    assign pp_31_24 = (select_e_31 & IN2[24] | select_2x_31 & IN2[23] | select_n2x_31 & (~ IN2[23]) | select_ne_31 & (~ IN2[24])  );
    wire logic pp_31_25;
    assign pp_31_25 = (select_e_31 & IN2[25] | select_2x_31 & IN2[24] | select_n2x_31 & (~ IN2[24]) | select_ne_31 & (~ IN2[25])  );
    wire logic pp_31_26;
    assign pp_31_26 = (select_e_31 & IN2[26] | select_2x_31 & IN2[25] | select_n2x_31 & (~ IN2[25]) | select_ne_31 & (~ IN2[26])  );
    wire logic pp_31_27;
    assign pp_31_27 = (select_e_31 & IN2[27] | select_2x_31 & IN2[26] | select_n2x_31 & (~ IN2[26]) | select_ne_31 & (~ IN2[27])  );
    wire logic pp_31_28;
    assign pp_31_28 = (select_e_31 & IN2[28] | select_2x_31 & IN2[27] | select_n2x_31 & (~ IN2[27]) | select_ne_31 & (~ IN2[28])  );
    wire logic pp_31_29;
    assign pp_31_29 = (select_e_31 & IN2[29] | select_2x_31 & IN2[28] | select_n2x_31 & (~ IN2[28]) | select_ne_31 & (~ IN2[29])  );
    wire logic pp_31_30;
    assign pp_31_30 = (select_e_31 & IN2[30] | select_2x_31 & IN2[29] | select_n2x_31 & (~ IN2[29]) | select_ne_31 & (~ IN2[30])  );
    wire logic pp_31_31;
    assign pp_31_31 = (select_e_31 & IN2[31] | select_2x_31 & IN2[30] | select_n2x_31 & (~ IN2[30]) | select_ne_31 & (~ IN2[31])  );
    wire logic pp_31_32;
    assign pp_31_32 = (select_e_31 & IN2[32] | select_2x_31 & IN2[31] | select_n2x_31 & (~ IN2[31]) | select_ne_31 & (~ IN2[32])  );
    wire logic pp_31_33;
    assign pp_31_33 = (select_e_31 & IN2[33] | select_2x_31 & IN2[32] | select_n2x_31 & (~ IN2[32]) | select_ne_31 & (~ IN2[33])  );
    wire logic pp_31_34;
    assign pp_31_34 = (select_e_31 & IN2[34] | select_2x_31 & IN2[33] | select_n2x_31 & (~ IN2[33]) | select_ne_31 & (~ IN2[34])  );
    wire logic pp_31_35;
    assign pp_31_35 = (select_e_31 & IN2[35] | select_2x_31 & IN2[34] | select_n2x_31 & (~ IN2[34]) | select_ne_31 & (~ IN2[35])  );
    wire logic pp_31_36;
    assign pp_31_36 = (select_e_31 & IN2[36] | select_2x_31 & IN2[35] | select_n2x_31 & (~ IN2[35]) | select_ne_31 & (~ IN2[36])  );
    wire logic pp_31_37;
    assign pp_31_37 = (select_e_31 & IN2[37] | select_2x_31 & IN2[36] | select_n2x_31 & (~ IN2[36]) | select_ne_31 & (~ IN2[37])  );
    wire logic pp_31_38;
    assign pp_31_38 = (select_e_31 & IN2[38] | select_2x_31 & IN2[37] | select_n2x_31 & (~ IN2[37]) | select_ne_31 & (~ IN2[38])  );
    wire logic pp_31_39;
    assign pp_31_39 = (select_e_31 & IN2[39] | select_2x_31 & IN2[38] | select_n2x_31 & (~ IN2[38]) | select_ne_31 & (~ IN2[39])  );
    wire logic pp_31_40;
    assign pp_31_40 = (select_e_31 & IN2[40] | select_2x_31 & IN2[39] | select_n2x_31 & (~ IN2[39]) | select_ne_31 & (~ IN2[40])  );
    wire logic pp_31_41;
    assign pp_31_41 = (select_e_31 & IN2[41] | select_2x_31 & IN2[40] | select_n2x_31 & (~ IN2[40]) | select_ne_31 & (~ IN2[41])  );
    wire logic pp_31_42;
    assign pp_31_42 = (select_e_31 & IN2[42] | select_2x_31 & IN2[41] | select_n2x_31 & (~ IN2[41]) | select_ne_31 & (~ IN2[42])  );
    wire logic pp_31_43;
    assign pp_31_43 = (select_e_31 & IN2[43] | select_2x_31 & IN2[42] | select_n2x_31 & (~ IN2[42]) | select_ne_31 & (~ IN2[43])  );
    wire logic pp_31_44;
    assign pp_31_44 = (select_e_31 & IN2[44] | select_2x_31 & IN2[43] | select_n2x_31 & (~ IN2[43]) | select_ne_31 & (~ IN2[44])  );
    wire logic pp_31_45;
    assign pp_31_45 = (select_e_31 & IN2[45] | select_2x_31 & IN2[44] | select_n2x_31 & (~ IN2[44]) | select_ne_31 & (~ IN2[45])  );
    wire logic pp_31_46;
    assign pp_31_46 = (select_e_31 & IN2[46] | select_2x_31 & IN2[45] | select_n2x_31 & (~ IN2[45]) | select_ne_31 & (~ IN2[46])  );
    wire logic pp_31_47;
    assign pp_31_47 = (select_e_31 & IN2[47] | select_2x_31 & IN2[46] | select_n2x_31 & (~ IN2[46]) | select_ne_31 & (~ IN2[47])  );
    wire logic pp_31_48;
    assign pp_31_48 = (select_e_31 & IN2[48] | select_2x_31 & IN2[47] | select_n2x_31 & (~ IN2[47]) | select_ne_31 & (~ IN2[48])  );
    wire logic pp_31_49;
    assign pp_31_49 = (select_e_31 & IN2[49] | select_2x_31 & IN2[48] | select_n2x_31 & (~ IN2[48]) | select_ne_31 & (~ IN2[49])  );
    wire logic pp_31_50;
    assign pp_31_50 = (select_e_31 & IN2[50] | select_2x_31 & IN2[49] | select_n2x_31 & (~ IN2[49]) | select_ne_31 & (~ IN2[50])  );
    wire logic pp_31_51;
    assign pp_31_51 = (select_e_31 & IN2[51] | select_2x_31 & IN2[50] | select_n2x_31 & (~ IN2[50]) | select_ne_31 & (~ IN2[51])  );
    wire logic pp_31_52;
    assign pp_31_52 = (select_e_31 & IN2[52] | select_2x_31 & IN2[51] | select_n2x_31 & (~ IN2[51]) | select_ne_31 & (~ IN2[52])  );
    wire logic pp_31_53;
    assign pp_31_53 = (select_e_31 & IN2[53] | select_2x_31 & IN2[52] | select_n2x_31 & (~ IN2[52]) | select_ne_31 & (~ IN2[53])  );
    wire logic pp_31_54;
    assign pp_31_54 = (select_e_31 & IN2[54] | select_2x_31 & IN2[53] | select_n2x_31 & (~ IN2[53]) | select_ne_31 & (~ IN2[54])  );
    wire logic pp_31_55;
    assign pp_31_55 = (select_e_31 & IN2[55] | select_2x_31 & IN2[54] | select_n2x_31 & (~ IN2[54]) | select_ne_31 & (~ IN2[55])  );
    wire logic pp_31_56;
    assign pp_31_56 = (select_e_31 & IN2[56] | select_2x_31 & IN2[55] | select_n2x_31 & (~ IN2[55]) | select_ne_31 & (~ IN2[56])  );
    wire logic pp_31_57;
    assign pp_31_57 = (select_e_31 & IN2[57] | select_2x_31 & IN2[56] | select_n2x_31 & (~ IN2[56]) | select_ne_31 & (~ IN2[57])  );
    wire logic pp_31_58;
    assign pp_31_58 = (select_e_31 & IN2[58] | select_2x_31 & IN2[57] | select_n2x_31 & (~ IN2[57]) | select_ne_31 & (~ IN2[58])  );
    wire logic pp_31_59;
    assign pp_31_59 = (select_e_31 & IN2[59] | select_2x_31 & IN2[58] | select_n2x_31 & (~ IN2[58]) | select_ne_31 & (~ IN2[59])  );
    wire logic pp_31_60;
    assign pp_31_60 = (select_e_31 & IN2[60] | select_2x_31 & IN2[59] | select_n2x_31 & (~ IN2[59]) | select_ne_31 & (~ IN2[60])  );
    wire logic pp_31_61;
    assign pp_31_61 = (select_e_31 & IN2[61] | select_2x_31 & IN2[60] | select_n2x_31 & (~ IN2[60]) | select_ne_31 & (~ IN2[61])  );
    wire logic pp_31_62;
    assign pp_31_62 = (select_e_31 & IN2[62] | select_2x_31 & IN2[61] | select_n2x_31 & (~ IN2[61]) | select_ne_31 & (~ IN2[62])  );
    wire logic pp_31_63;
    assign pp_31_63 = (select_e_31 & IN2[63] | select_2x_31 & IN2[62] | select_n2x_31 & (~ IN2[62]) | select_ne_31 & (~ IN2[63])  );
    wire logic pp_31_64;
    assign pp_31_64 = (select_e_31 & IN2[63] | select_2x_31 & IN2[63] | select_n2x_31 & (~ IN2[63]) | select_ne_31 & (~ IN2[63])  );
    wire logic pp_31_65;
    assign pp_31_65 = ~ (select_e_31 & IN2[63] | select_2x_31 & IN2[63] | select_n2x_31 & (~ IN2[63]) | select_ne_31 & (~ IN2[63])  );
    assign tcomp31 = select_ne_31 | select_n2x_31;
    
// Creating Summation Tree 

    logic s0 ,c0;
    ha ha0 (pp_0_54, pp_1_52, s0, c0);
    logic s1 ,c1;
    ha ha1 (pp_0_55, pp_1_53, s1, c1);
    logic s2 ,c2; 
    fa fa2 (pp_0_56, pp_1_54, pp_2_52, s2, c2);
    logic s3 ,c3;
    ha ha3 (pp_3_50, pp_4_48, s3, c3);
    logic s4 ,c4; 
    fa fa4 (pp_0_57, pp_1_55, pp_2_53, s4, c4);
    logic s5 ,c5;
    ha ha5 (pp_3_51, pp_4_49, s5, c5);
    logic s6 ,c6; 
    fa fa6 (pp_0_58, pp_1_56, pp_2_54, s6, c6);
    logic s7 ,c7; 
    fa fa7 (pp_3_52, pp_4_50, pp_5_48, s7, c7);
    logic s8 ,c8;
    ha ha8 (pp_6_46, pp_7_44, s8, c8);
    logic s9 ,c9; 
    fa fa9 (pp_0_59, pp_1_57, pp_2_55, s9, c9);
    logic s10 ,c10; 
    fa fa10 (pp_3_53, pp_4_51, pp_5_49, s10, c10);
    logic s11 ,c11;
    ha ha11 (pp_6_47, pp_7_45, s11, c11);
    logic s12 ,c12; 
    fa fa12 (pp_0_60, pp_1_58, pp_2_56, s12, c12);
    logic s13 ,c13; 
    fa fa13 (pp_3_54, pp_4_52, pp_5_50, s13, c13);
    logic s14 ,c14; 
    fa fa14 (pp_6_48, pp_7_46, pp_8_44, s14, c14);
    logic s15 ,c15;
    ha ha15 (pp_9_42, pp_10_40, s15, c15);
    logic s16 ,c16; 
    fa fa16 (pp_0_61, pp_1_59, pp_2_57, s16, c16);
    logic s17 ,c17; 
    fa fa17 (pp_3_55, pp_4_53, pp_5_51, s17, c17);
    logic s18 ,c18; 
    fa fa18 (pp_6_49, pp_7_47, pp_8_45, s18, c18);
    logic s19 ,c19;
    ha ha19 (pp_9_43, pp_10_41, s19, c19);
    logic s20 ,c20; 
    fa fa20 (pp_0_62, pp_1_60, pp_2_58, s20, c20);
    logic s21 ,c21; 
    fa fa21 (pp_3_56, pp_4_54, pp_5_52, s21, c21);
    logic s22 ,c22; 
    fa fa22 (pp_6_50, pp_7_48, pp_8_46, s22, c22);
    logic s23 ,c23; 
    fa fa23 (pp_9_44, pp_10_42, pp_11_40, s23, c23);
    logic s24 ,c24;
    ha ha24 (pp_12_38, pp_13_36, s24, c24);
    logic s25 ,c25; 
    fa fa25 (pp_0_63, pp_1_61, pp_2_59, s25, c25);
    logic s26 ,c26; 
    fa fa26 (pp_3_57, pp_4_55, pp_5_53, s26, c26);
    logic s27 ,c27; 
    fa fa27 (pp_6_51, pp_7_49, pp_8_47, s27, c27);
    logic s28 ,c28; 
    fa fa28 (pp_9_45, pp_10_43, pp_11_41, s28, c28);
    logic s29 ,c29;
    ha ha29 (pp_12_39, pp_13_37, s29, c29);
    logic s30 ,c30; 
    fa fa30 (pp_0_64, pp_1_62, pp_2_60, s30, c30);
    logic s31 ,c31; 
    fa fa31 (pp_3_58, pp_4_56, pp_5_54, s31, c31);
    logic s32 ,c32; 
    fa fa32 (pp_6_52, pp_7_50, pp_8_48, s32, c32);
    logic s33 ,c33; 
    fa fa33 (pp_9_46, pp_10_44, pp_11_42, s33, c33);
    logic s34 ,c34;
    ha ha34 (pp_12_40, pp_13_38, s34, c34);
    logic s35 ,c35; 
    fa fa35 (pp_0_65, pp_1_63, pp_2_61, s35, c35);
    logic s36 ,c36; 
    fa fa36 (pp_3_59, pp_4_57, pp_5_55, s36, c36);
    logic s37 ,c37; 
    fa fa37 (pp_6_53, pp_7_51, pp_8_49, s37, c37);
    logic s38 ,c38; 
    fa fa38 (pp_9_47, pp_10_45, pp_11_43, s38, c38);
    logic s39 ,c39; 
    fa fa39 (pp_12_41, pp_13_39, pp_14_37, s39, c39);
    logic s40 ,c40; 
    fa fa40 (const1, pp_1_64, pp_2_62, s40, c40);
    logic s41 ,c41; 
    fa fa41 (pp_3_60, pp_4_58, pp_5_56, s41, c41);
    logic s42 ,c42; 
    fa fa42 (pp_6_54, pp_7_52, pp_8_50, s42, c42);
    logic s43 ,c43; 
    fa fa43 (pp_9_48, pp_10_46, pp_11_44, s43, c43);
    logic s44 ,c44;
    ha ha44 (pp_12_42, pp_13_40, s44, c44);
    logic s45 ,c45; 
    fa fa45 (pp_1_65, pp_2_63, pp_3_61, s45, c45);
    logic s46 ,c46; 
    fa fa46 (pp_4_59, pp_5_57, pp_6_55, s46, c46);
    logic s47 ,c47; 
    fa fa47 (pp_7_53, pp_8_51, pp_9_49, s47, c47);
    logic s48 ,c48; 
    fa fa48 (pp_10_47, pp_11_45, pp_12_43, s48, c48);
    logic s49 ,c49; 
    fa fa49 (const1, pp_2_64, pp_3_62, s49, c49);
    logic s50 ,c50; 
    fa fa50 (pp_4_60, pp_5_58, pp_6_56, s50, c50);
    logic s51 ,c51; 
    fa fa51 (pp_7_54, pp_8_52, pp_9_50, s51, c51);
    logic s52 ,c52;
    ha ha52 (pp_10_48, pp_11_46, s52, c52);
    logic s53 ,c53; 
    fa fa53 (pp_2_65, pp_3_63, pp_4_61, s53, c53);
    logic s54 ,c54; 
    fa fa54 (pp_5_59, pp_6_57, pp_7_55, s54, c54);
    logic s55 ,c55; 
    fa fa55 (pp_8_53, pp_9_51, pp_10_49, s55, c55);
    logic s56 ,c56; 
    fa fa56 (const1, pp_3_64, pp_4_62, s56, c56);
    logic s57 ,c57; 
    fa fa57 (pp_5_60, pp_6_58, pp_7_56, s57, c57);
    logic s58 ,c58;
    ha ha58 (pp_8_54, pp_9_52, s58, c58);
    logic s59 ,c59; 
    fa fa59 (pp_3_65, pp_4_63, pp_5_61, s59, c59);
    logic s60 ,c60; 
    fa fa60 (pp_6_59, pp_7_57, pp_8_55, s60, c60);
    logic s61 ,c61; 
    fa fa61 (const1, pp_4_64, pp_5_62, s61, c61);
    logic s62 ,c62;
    ha ha62 (pp_6_60, pp_7_58, s62, c62);
    logic s63 ,c63; 
    fa fa63 (pp_4_65, pp_5_63, pp_6_61, s63, c63);
    logic s64 ,c64;
    ha ha64 (const1, pp_5_64, s64, c64);
    logic s65 ,c65;
    ha ha65 (pp_0_36, pp_1_34, s65, c65);
    logic s66 ,c66;
    ha ha66 (pp_0_37, pp_1_35, s66, c66);
    logic s67 ,c67; 
    fa fa67 (pp_0_38, pp_1_36, pp_2_34, s67, c67);
    logic s68 ,c68;
    ha ha68 (pp_3_32, pp_4_30, s68, c68);
    logic s69 ,c69; 
    fa fa69 (pp_0_39, pp_1_37, pp_2_35, s69, c69);
    logic s70 ,c70;
    ha ha70 (pp_3_33, pp_4_31, s70, c70);
    logic s71 ,c71; 
    fa fa71 (pp_0_40, pp_1_38, pp_2_36, s71, c71);
    logic s72 ,c72; 
    fa fa72 (pp_3_34, pp_4_32, pp_5_30, s72, c72);
    logic s73 ,c73;
    ha ha73 (pp_6_28, pp_7_26, s73, c73);
    logic s74 ,c74; 
    fa fa74 (pp_0_41, pp_1_39, pp_2_37, s74, c74);
    logic s75 ,c75; 
    fa fa75 (pp_3_35, pp_4_33, pp_5_31, s75, c75);
    logic s76 ,c76;
    ha ha76 (pp_6_29, pp_7_27, s76, c76);
    logic s77 ,c77; 
    fa fa77 (pp_0_42, pp_1_40, pp_2_38, s77, c77);
    logic s78 ,c78; 
    fa fa78 (pp_3_36, pp_4_34, pp_5_32, s78, c78);
    logic s79 ,c79; 
    fa fa79 (pp_6_30, pp_7_28, pp_8_26, s79, c79);
    logic s80 ,c80;
    ha ha80 (pp_9_24, pp_10_22, s80, c80);
    logic s81 ,c81; 
    fa fa81 (pp_0_43, pp_1_41, pp_2_39, s81, c81);
    logic s82 ,c82; 
    fa fa82 (pp_3_37, pp_4_35, pp_5_33, s82, c82);
    logic s83 ,c83; 
    fa fa83 (pp_6_31, pp_7_29, pp_8_27, s83, c83);
    logic s84 ,c84;
    ha ha84 (pp_9_25, pp_10_23, s84, c84);
    logic s85 ,c85; 
    fa fa85 (pp_0_44, pp_1_42, pp_2_40, s85, c85);
    logic s86 ,c86; 
    fa fa86 (pp_3_38, pp_4_36, pp_5_34, s86, c86);
    logic s87 ,c87; 
    fa fa87 (pp_6_32, pp_7_30, pp_8_28, s87, c87);
    logic s88 ,c88; 
    fa fa88 (pp_9_26, pp_10_24, pp_11_22, s88, c88);
    logic s89 ,c89;
    ha ha89 (pp_12_20, pp_13_18, s89, c89);
    logic s90 ,c90; 
    fa fa90 (pp_0_45, pp_1_43, pp_2_41, s90, c90);
    logic s91 ,c91; 
    fa fa91 (pp_3_39, pp_4_37, pp_5_35, s91, c91);
    logic s92 ,c92; 
    fa fa92 (pp_6_33, pp_7_31, pp_8_29, s92, c92);
    logic s93 ,c93; 
    fa fa93 (pp_9_27, pp_10_25, pp_11_23, s93, c93);
    logic s94 ,c94;
    ha ha94 (pp_12_21, pp_13_19, s94, c94);
    logic s95 ,c95; 
    fa fa95 (pp_0_46, pp_1_44, pp_2_42, s95, c95);
    logic s96 ,c96; 
    fa fa96 (pp_3_40, pp_4_38, pp_5_36, s96, c96);
    logic s97 ,c97; 
    fa fa97 (pp_6_34, pp_7_32, pp_8_30, s97, c97);
    logic s98 ,c98; 
    fa fa98 (pp_9_28, pp_10_26, pp_11_24, s98, c98);
    logic s99 ,c99; 
    fa fa99 (pp_12_22, pp_13_20, pp_14_18, s99, c99);
    logic s100 ,c100;
    ha ha100 (pp_15_16, pp_16_14, s100, c100);
    logic s101 ,c101; 
    fa fa101 (pp_0_47, pp_1_45, pp_2_43, s101, c101);
    logic s102 ,c102; 
    fa fa102 (pp_3_41, pp_4_39, pp_5_37, s102, c102);
    logic s103 ,c103; 
    fa fa103 (pp_6_35, pp_7_33, pp_8_31, s103, c103);
    logic s104 ,c104; 
    fa fa104 (pp_9_29, pp_10_27, pp_11_25, s104, c104);
    logic s105 ,c105; 
    fa fa105 (pp_12_23, pp_13_21, pp_14_19, s105, c105);
    logic s106 ,c106;
    ha ha106 (pp_15_17, pp_16_15, s106, c106);
    logic s107 ,c107; 
    fa fa107 (pp_0_48, pp_1_46, pp_2_44, s107, c107);
    logic s108 ,c108; 
    fa fa108 (pp_3_42, pp_4_40, pp_5_38, s108, c108);
    logic s109 ,c109; 
    fa fa109 (pp_6_36, pp_7_34, pp_8_32, s109, c109);
    logic s110 ,c110; 
    fa fa110 (pp_9_30, pp_10_28, pp_11_26, s110, c110);
    logic s111 ,c111; 
    fa fa111 (pp_12_24, pp_13_22, pp_14_20, s111, c111);
    logic s112 ,c112; 
    fa fa112 (pp_15_18, pp_16_16, pp_17_14, s112, c112);
    logic s113 ,c113;
    ha ha113 (pp_18_12, pp_19_10, s113, c113);
    logic s114 ,c114; 
    fa fa114 (pp_0_49, pp_1_47, pp_2_45, s114, c114);
    logic s115 ,c115; 
    fa fa115 (pp_3_43, pp_4_41, pp_5_39, s115, c115);
    logic s116 ,c116; 
    fa fa116 (pp_6_37, pp_7_35, pp_8_33, s116, c116);
    logic s117 ,c117; 
    fa fa117 (pp_9_31, pp_10_29, pp_11_27, s117, c117);
    logic s118 ,c118; 
    fa fa118 (pp_12_25, pp_13_23, pp_14_21, s118, c118);
    logic s119 ,c119; 
    fa fa119 (pp_15_19, pp_16_17, pp_17_15, s119, c119);
    logic s120 ,c120;
    ha ha120 (pp_18_13, pp_19_11, s120, c120);
    logic s121 ,c121; 
    fa fa121 (pp_0_50, pp_1_48, pp_2_46, s121, c121);
    logic s122 ,c122; 
    fa fa122 (pp_3_44, pp_4_42, pp_5_40, s122, c122);
    logic s123 ,c123; 
    fa fa123 (pp_6_38, pp_7_36, pp_8_34, s123, c123);
    logic s124 ,c124; 
    fa fa124 (pp_9_32, pp_10_30, pp_11_28, s124, c124);
    logic s125 ,c125; 
    fa fa125 (pp_12_26, pp_13_24, pp_14_22, s125, c125);
    logic s126 ,c126; 
    fa fa126 (pp_15_20, pp_16_18, pp_17_16, s126, c126);
    logic s127 ,c127; 
    fa fa127 (pp_18_14, pp_19_12, pp_20_10, s127, c127);
    logic s128 ,c128;
    ha ha128 (pp_21_8, pp_22_6, s128, c128);
    logic s129 ,c129; 
    fa fa129 (pp_0_51, pp_1_49, pp_2_47, s129, c129);
    logic s130 ,c130; 
    fa fa130 (pp_3_45, pp_4_43, pp_5_41, s130, c130);
    logic s131 ,c131; 
    fa fa131 (pp_6_39, pp_7_37, pp_8_35, s131, c131);
    logic s132 ,c132; 
    fa fa132 (pp_9_33, pp_10_31, pp_11_29, s132, c132);
    logic s133 ,c133; 
    fa fa133 (pp_12_27, pp_13_25, pp_14_23, s133, c133);
    logic s134 ,c134; 
    fa fa134 (pp_15_21, pp_16_19, pp_17_17, s134, c134);
    logic s135 ,c135; 
    fa fa135 (pp_18_15, pp_19_13, pp_20_11, s135, c135);
    logic s136 ,c136;
    ha ha136 (pp_21_9, pp_22_7, s136, c136);
    logic s137 ,c137; 
    fa fa137 (pp_0_52, pp_1_50, pp_2_48, s137, c137);
    logic s138 ,c138; 
    fa fa138 (pp_3_46, pp_4_44, pp_5_42, s138, c138);
    logic s139 ,c139; 
    fa fa139 (pp_6_40, pp_7_38, pp_8_36, s139, c139);
    logic s140 ,c140; 
    fa fa140 (pp_9_34, pp_10_32, pp_11_30, s140, c140);
    logic s141 ,c141; 
    fa fa141 (pp_12_28, pp_13_26, pp_14_24, s141, c141);
    logic s142 ,c142; 
    fa fa142 (pp_15_22, pp_16_20, pp_17_18, s142, c142);
    logic s143 ,c143; 
    fa fa143 (pp_18_16, pp_19_14, pp_20_12, s143, c143);
    logic s144 ,c144; 
    fa fa144 (pp_21_10, pp_22_8, pp_23_6, s144, c144);
    logic s145 ,c145;
    ha ha145 (pp_24_4, pp_25_2, s145, c145);
    logic s146 ,c146; 
    fa fa146 (pp_0_53, pp_1_51, pp_2_49, s146, c146);
    logic s147 ,c147; 
    fa fa147 (pp_3_47, pp_4_45, pp_5_43, s147, c147);
    logic s148 ,c148; 
    fa fa148 (pp_6_41, pp_7_39, pp_8_37, s148, c148);
    logic s149 ,c149; 
    fa fa149 (pp_9_35, pp_10_33, pp_11_31, s149, c149);
    logic s150 ,c150; 
    fa fa150 (pp_12_29, pp_13_27, pp_14_25, s150, c150);
    logic s151 ,c151; 
    fa fa151 (pp_15_23, pp_16_21, pp_17_19, s151, c151);
    logic s152 ,c152; 
    fa fa152 (pp_18_17, pp_19_15, pp_20_13, s152, c152);
    logic s153 ,c153; 
    fa fa153 (pp_21_11, pp_22_9, pp_23_7, s153, c153);
    logic s154 ,c154;
    ha ha154 (pp_24_5, pp_25_3, s154, c154);
    logic s155 ,c155; 
    fa fa155 (pp_2_50, pp_3_48, pp_4_46, s155, c155);
    logic s156 ,c156; 
    fa fa156 (pp_5_44, pp_6_42, pp_7_40, s156, c156);
    logic s157 ,c157; 
    fa fa157 (pp_8_38, pp_9_36, pp_10_34, s157, c157);
    logic s158 ,c158; 
    fa fa158 (pp_11_32, pp_12_30, pp_13_28, s158, c158);
    logic s159 ,c159; 
    fa fa159 (pp_14_26, pp_15_24, pp_16_22, s159, c159);
    logic s160 ,c160; 
    fa fa160 (pp_17_20, pp_18_18, pp_19_16, s160, c160);
    logic s161 ,c161; 
    fa fa161 (pp_20_14, pp_21_12, pp_22_10, s161, c161);
    logic s162 ,c162; 
    fa fa162 (pp_23_8, pp_24_6, pp_25_4, s162, c162);
    logic s163 ,c163; 
    fa fa163 (pp_26_2, pp_27_0, tcomp27, s163, c163);
    logic s164 ,c164; 
    fa fa164 (pp_2_51, pp_3_49, pp_4_47, s164, c164);
    logic s165 ,c165; 
    fa fa165 (pp_5_45, pp_6_43, pp_7_41, s165, c165);
    logic s166 ,c166; 
    fa fa166 (pp_8_39, pp_9_37, pp_10_35, s166, c166);
    logic s167 ,c167; 
    fa fa167 (pp_11_33, pp_12_31, pp_13_29, s167, c167);
    logic s168 ,c168; 
    fa fa168 (pp_14_27, pp_15_25, pp_16_23, s168, c168);
    logic s169 ,c169; 
    fa fa169 (pp_17_21, pp_18_19, pp_19_17, s169, c169);
    logic s170 ,c170; 
    fa fa170 (pp_20_15, pp_21_13, pp_22_11, s170, c170);
    logic s171 ,c171; 
    fa fa171 (pp_23_9, pp_24_7, pp_25_5, s171, c171);
    logic s172 ,c172; 
    fa fa172 (pp_26_3, pp_27_1, c0, s172, c172);
    logic s173 ,c173; 
    fa fa173 (pp_5_46, pp_6_44, pp_7_42, s173, c173);
    logic s174 ,c174; 
    fa fa174 (pp_8_40, pp_9_38, pp_10_36, s174, c174);
    logic s175 ,c175; 
    fa fa175 (pp_11_34, pp_12_32, pp_13_30, s175, c175);
    logic s176 ,c176; 
    fa fa176 (pp_14_28, pp_15_26, pp_16_24, s176, c176);
    logic s177 ,c177; 
    fa fa177 (pp_17_22, pp_18_20, pp_19_18, s177, c177);
    logic s178 ,c178; 
    fa fa178 (pp_20_16, pp_21_14, pp_22_12, s178, c178);
    logic s179 ,c179; 
    fa fa179 (pp_23_10, pp_24_8, pp_25_6, s179, c179);
    logic s180 ,c180; 
    fa fa180 (pp_26_4, pp_27_2, pp_28_0, s180, c180);
    logic s181 ,c181; 
    fa fa181 (tcomp28, c1, s2, s181, c181);
    logic s182 ,c182; 
    fa fa182 (pp_5_47, pp_6_45, pp_7_43, s182, c182);
    logic s183 ,c183; 
    fa fa183 (pp_8_41, pp_9_39, pp_10_37, s183, c183);
    logic s184 ,c184; 
    fa fa184 (pp_11_35, pp_12_33, pp_13_31, s184, c184);
    logic s185 ,c185; 
    fa fa185 (pp_14_29, pp_15_27, pp_16_25, s185, c185);
    logic s186 ,c186; 
    fa fa186 (pp_17_23, pp_18_21, pp_19_19, s186, c186);
    logic s187 ,c187; 
    fa fa187 (pp_20_17, pp_21_15, pp_22_13, s187, c187);
    logic s188 ,c188; 
    fa fa188 (pp_23_11, pp_24_9, pp_25_7, s188, c188);
    logic s189 ,c189; 
    fa fa189 (pp_26_5, pp_27_3, pp_28_1, s189, c189);
    logic s190 ,c190; 
    fa fa190 (c2, c3, s4, s190, c190);
    logic s191 ,c191; 
    fa fa191 (pp_8_42, pp_9_40, pp_10_38, s191, c191);
    logic s192 ,c192; 
    fa fa192 (pp_11_36, pp_12_34, pp_13_32, s192, c192);
    logic s193 ,c193; 
    fa fa193 (pp_14_30, pp_15_28, pp_16_26, s193, c193);
    logic s194 ,c194; 
    fa fa194 (pp_17_24, pp_18_22, pp_19_20, s194, c194);
    logic s195 ,c195; 
    fa fa195 (pp_20_18, pp_21_16, pp_22_14, s195, c195);
    logic s196 ,c196; 
    fa fa196 (pp_23_12, pp_24_10, pp_25_8, s196, c196);
    logic s197 ,c197; 
    fa fa197 (pp_26_6, pp_27_4, pp_28_2, s197, c197);
    logic s198 ,c198; 
    fa fa198 (pp_29_0, tcomp29, c4, s198, c198);
    logic s199 ,c199; 
    fa fa199 (c5, s6, s7, s199, c199);
    logic s200 ,c200; 
    fa fa200 (pp_8_43, pp_9_41, pp_10_39, s200, c200);
    logic s201 ,c201; 
    fa fa201 (pp_11_37, pp_12_35, pp_13_33, s201, c201);
    logic s202 ,c202; 
    fa fa202 (pp_14_31, pp_15_29, pp_16_27, s202, c202);
    logic s203 ,c203; 
    fa fa203 (pp_17_25, pp_18_23, pp_19_21, s203, c203);
    logic s204 ,c204; 
    fa fa204 (pp_20_19, pp_21_17, pp_22_15, s204, c204);
    logic s205 ,c205; 
    fa fa205 (pp_23_13, pp_24_11, pp_25_9, s205, c205);
    logic s206 ,c206; 
    fa fa206 (pp_26_7, pp_27_5, pp_28_3, s206, c206);
    logic s207 ,c207; 
    fa fa207 (pp_29_1, c6, c7, s207, c207);
    logic s208 ,c208; 
    fa fa208 (c8, s9, s10, s208, c208);
    logic s209 ,c209; 
    fa fa209 (pp_11_38, pp_12_36, pp_13_34, s209, c209);
    logic s210 ,c210; 
    fa fa210 (pp_14_32, pp_15_30, pp_16_28, s210, c210);
    logic s211 ,c211; 
    fa fa211 (pp_17_26, pp_18_24, pp_19_22, s211, c211);
    logic s212 ,c212; 
    fa fa212 (pp_20_20, pp_21_18, pp_22_16, s212, c212);
    logic s213 ,c213; 
    fa fa213 (pp_23_14, pp_24_12, pp_25_10, s213, c213);
    logic s214 ,c214; 
    fa fa214 (pp_26_8, pp_27_6, pp_28_4, s214, c214);
    logic s215 ,c215; 
    fa fa215 (pp_29_2, pp_30_0, tcomp30, s215, c215);
    logic s216 ,c216; 
    fa fa216 (c9, c10, c11, s216, c216);
    logic s217 ,c217; 
    fa fa217 (s12, s13, s14, s217, c217);
    logic s218 ,c218; 
    fa fa218 (pp_11_39, pp_12_37, pp_13_35, s218, c218);
    logic s219 ,c219; 
    fa fa219 (pp_14_33, pp_15_31, pp_16_29, s219, c219);
    logic s220 ,c220; 
    fa fa220 (pp_17_27, pp_18_25, pp_19_23, s220, c220);
    logic s221 ,c221; 
    fa fa221 (pp_20_21, pp_21_19, pp_22_17, s221, c221);
    logic s222 ,c222; 
    fa fa222 (pp_23_15, pp_24_13, pp_25_11, s222, c222);
    logic s223 ,c223; 
    fa fa223 (pp_26_9, pp_27_7, pp_28_5, s223, c223);
    logic s224 ,c224; 
    fa fa224 (pp_29_3, pp_30_1, c12, s224, c224);
    logic s225 ,c225; 
    fa fa225 (c13, c14, c15, s225, c225);
    logic s226 ,c226; 
    fa fa226 (s16, s17, s18, s226, c226);
    logic s227 ,c227; 
    fa fa227 (pp_14_34, pp_15_32, pp_16_30, s227, c227);
    logic s228 ,c228; 
    fa fa228 (pp_17_28, pp_18_26, pp_19_24, s228, c228);
    logic s229 ,c229; 
    fa fa229 (pp_20_22, pp_21_20, pp_22_18, s229, c229);
    logic s230 ,c230; 
    fa fa230 (pp_23_16, pp_24_14, pp_25_12, s230, c230);
    logic s231 ,c231; 
    fa fa231 (pp_26_10, pp_27_8, pp_28_6, s231, c231);
    logic s232 ,c232; 
    fa fa232 (pp_29_4, pp_30_2, pp_31_0, s232, c232);
    logic s233 ,c233; 
    fa fa233 (tcomp31, c16, c17, s233, c233);
    logic s234 ,c234; 
    fa fa234 (c18, c19, s20, s234, c234);
    logic s235 ,c235; 
    fa fa235 (s21, s22, s23, s235, c235);
    logic s236 ,c236; 
    fa fa236 (pp_14_35, pp_15_33, pp_16_31, s236, c236);
    logic s237 ,c237; 
    fa fa237 (pp_17_29, pp_18_27, pp_19_25, s237, c237);
    logic s238 ,c238; 
    fa fa238 (pp_20_23, pp_21_21, pp_22_19, s238, c238);
    logic s239 ,c239; 
    fa fa239 (pp_23_17, pp_24_15, pp_25_13, s239, c239);
    logic s240 ,c240; 
    fa fa240 (pp_26_11, pp_27_9, pp_28_7, s240, c240);
    logic s241 ,c241; 
    fa fa241 (pp_29_5, pp_30_3, pp_31_1, s241, c241);
    logic s242 ,c242; 
    fa fa242 (c20, c21, c22, s242, c242);
    logic s243 ,c243; 
    fa fa243 (c23, c24, s25, s243, c243);
    logic s244 ,c244; 
    fa fa244 (s26, s27, s28, s244, c244);
    logic s245 ,c245; 
    fa fa245 (pp_14_36, pp_15_34, pp_16_32, s245, c245);
    logic s246 ,c246; 
    fa fa246 (pp_17_30, pp_18_28, pp_19_26, s246, c246);
    logic s247 ,c247; 
    fa fa247 (pp_20_24, pp_21_22, pp_22_20, s247, c247);
    logic s248 ,c248; 
    fa fa248 (pp_23_18, pp_24_16, pp_25_14, s248, c248);
    logic s249 ,c249; 
    fa fa249 (pp_26_12, pp_27_10, pp_28_8, s249, c249);
    logic s250 ,c250; 
    fa fa250 (pp_29_6, pp_30_4, pp_31_2, s250, c250);
    logic s251 ,c251; 
    fa fa251 (c25, c26, c27, s251, c251);
    logic s252 ,c252; 
    fa fa252 (c28, c29, s30, s252, c252);
    logic s253 ,c253; 
    fa fa253 (s31, s32, s33, s253, c253);
    logic s254 ,c254; 
    fa fa254 (pp_15_35, pp_16_33, pp_17_31, s254, c254);
    logic s255 ,c255; 
    fa fa255 (pp_18_29, pp_19_27, pp_20_25, s255, c255);
    logic s256 ,c256; 
    fa fa256 (pp_21_23, pp_22_21, pp_23_19, s256, c256);
    logic s257 ,c257; 
    fa fa257 (pp_24_17, pp_25_15, pp_26_13, s257, c257);
    logic s258 ,c258; 
    fa fa258 (pp_27_11, pp_28_9, pp_29_7, s258, c258);
    logic s259 ,c259; 
    fa fa259 (pp_30_5, pp_31_3, const1, s259, c259);
    logic s260 ,c260; 
    fa fa260 (c30, c31, c32, s260, c260);
    logic s261 ,c261; 
    fa fa261 (c33, c34, s35, s261, c261);
    logic s262 ,c262; 
    fa fa262 (s36, s37, s38, s262, c262);
    logic s263 ,c263; 
    fa fa263 (pp_14_38, pp_15_36, pp_16_34, s263, c263);
    logic s264 ,c264; 
    fa fa264 (pp_17_32, pp_18_30, pp_19_28, s264, c264);
    logic s265 ,c265; 
    fa fa265 (pp_20_26, pp_21_24, pp_22_22, s265, c265);
    logic s266 ,c266; 
    fa fa266 (pp_23_20, pp_24_18, pp_25_16, s266, c266);
    logic s267 ,c267; 
    fa fa267 (pp_26_14, pp_27_12, pp_28_10, s267, c267);
    logic s268 ,c268; 
    fa fa268 (pp_29_8, pp_30_6, pp_31_4, s268, c268);
    logic s269 ,c269; 
    fa fa269 (c35, c36, c37, s269, c269);
    logic s270 ,c270; 
    fa fa270 (c38, c39, s40, s270, c270);
    logic s271 ,c271; 
    fa fa271 (s41, s42, s43, s271, c271);
    logic s272 ,c272; 
    fa fa272 (pp_13_41, pp_14_39, pp_15_37, s272, c272);
    logic s273 ,c273; 
    fa fa273 (pp_16_35, pp_17_33, pp_18_31, s273, c273);
    logic s274 ,c274; 
    fa fa274 (pp_19_29, pp_20_27, pp_21_25, s274, c274);
    logic s275 ,c275; 
    fa fa275 (pp_22_23, pp_23_21, pp_24_19, s275, c275);
    logic s276 ,c276; 
    fa fa276 (pp_25_17, pp_26_15, pp_27_13, s276, c276);
    logic s277 ,c277; 
    fa fa277 (pp_28_11, pp_29_9, pp_30_7, s277, c277);
    logic s278 ,c278; 
    fa fa278 (pp_31_5, c40, c41, s278, c278);
    logic s279 ,c279; 
    fa fa279 (c42, c43, c44, s279, c279);
    logic s280 ,c280; 
    fa fa280 (s45, s46, s47, s280, c280);
    logic s281 ,c281; 
    fa fa281 (pp_12_44, pp_13_42, pp_14_40, s281, c281);
    logic s282 ,c282; 
    fa fa282 (pp_15_38, pp_16_36, pp_17_34, s282, c282);
    logic s283 ,c283; 
    fa fa283 (pp_18_32, pp_19_30, pp_20_28, s283, c283);
    logic s284 ,c284; 
    fa fa284 (pp_21_26, pp_22_24, pp_23_22, s284, c284);
    logic s285 ,c285; 
    fa fa285 (pp_24_20, pp_25_18, pp_26_16, s285, c285);
    logic s286 ,c286; 
    fa fa286 (pp_27_14, pp_28_12, pp_29_10, s286, c286);
    logic s287 ,c287; 
    fa fa287 (pp_30_8, pp_31_6, c45, s287, c287);
    logic s288 ,c288; 
    fa fa288 (c46, c47, c48, s288, c288);
    logic s289 ,c289; 
    fa fa289 (s49, s50, s51, s289, c289);
    logic s290 ,c290; 
    fa fa290 (pp_11_47, pp_12_45, pp_13_43, s290, c290);
    logic s291 ,c291; 
    fa fa291 (pp_14_41, pp_15_39, pp_16_37, s291, c291);
    logic s292 ,c292; 
    fa fa292 (pp_17_35, pp_18_33, pp_19_31, s292, c292);
    logic s293 ,c293; 
    fa fa293 (pp_20_29, pp_21_27, pp_22_25, s293, c293);
    logic s294 ,c294; 
    fa fa294 (pp_23_23, pp_24_21, pp_25_19, s294, c294);
    logic s295 ,c295; 
    fa fa295 (pp_26_17, pp_27_15, pp_28_13, s295, c295);
    logic s296 ,c296; 
    fa fa296 (pp_29_11, pp_30_9, pp_31_7, s296, c296);
    logic s297 ,c297; 
    fa fa297 (c49, c50, c51, s297, c297);
    logic s298 ,c298; 
    fa fa298 (c52, s53, s54, s298, c298);
    logic s299 ,c299; 
    fa fa299 (pp_10_50, pp_11_48, pp_12_46, s299, c299);
    logic s300 ,c300; 
    fa fa300 (pp_13_44, pp_14_42, pp_15_40, s300, c300);
    logic s301 ,c301; 
    fa fa301 (pp_16_38, pp_17_36, pp_18_34, s301, c301);
    logic s302 ,c302; 
    fa fa302 (pp_19_32, pp_20_30, pp_21_28, s302, c302);
    logic s303 ,c303; 
    fa fa303 (pp_22_26, pp_23_24, pp_24_22, s303, c303);
    logic s304 ,c304; 
    fa fa304 (pp_25_20, pp_26_18, pp_27_16, s304, c304);
    logic s305 ,c305; 
    fa fa305 (pp_28_14, pp_29_12, pp_30_10, s305, c305);
    logic s306 ,c306; 
    fa fa306 (pp_31_8, c53, c54, s306, c306);
    logic s307 ,c307; 
    fa fa307 (c55, s56, s57, s307, c307);
    logic s308 ,c308; 
    fa fa308 (pp_9_53, pp_10_51, pp_11_49, s308, c308);
    logic s309 ,c309; 
    fa fa309 (pp_12_47, pp_13_45, pp_14_43, s309, c309);
    logic s310 ,c310; 
    fa fa310 (pp_15_41, pp_16_39, pp_17_37, s310, c310);
    logic s311 ,c311; 
    fa fa311 (pp_18_35, pp_19_33, pp_20_31, s311, c311);
    logic s312 ,c312; 
    fa fa312 (pp_21_29, pp_22_27, pp_23_25, s312, c312);
    logic s313 ,c313; 
    fa fa313 (pp_24_23, pp_25_21, pp_26_19, s313, c313);
    logic s314 ,c314; 
    fa fa314 (pp_27_17, pp_28_15, pp_29_13, s314, c314);
    logic s315 ,c315; 
    fa fa315 (pp_30_11, pp_31_9, c56, s315, c315);
    logic s316 ,c316; 
    fa fa316 (c57, c58, s59, s316, c316);
    logic s317 ,c317; 
    fa fa317 (pp_8_56, pp_9_54, pp_10_52, s317, c317);
    logic s318 ,c318; 
    fa fa318 (pp_11_50, pp_12_48, pp_13_46, s318, c318);
    logic s319 ,c319; 
    fa fa319 (pp_14_44, pp_15_42, pp_16_40, s319, c319);
    logic s320 ,c320; 
    fa fa320 (pp_17_38, pp_18_36, pp_19_34, s320, c320);
    logic s321 ,c321; 
    fa fa321 (pp_20_32, pp_21_30, pp_22_28, s321, c321);
    logic s322 ,c322; 
    fa fa322 (pp_23_26, pp_24_24, pp_25_22, s322, c322);
    logic s323 ,c323; 
    fa fa323 (pp_26_20, pp_27_18, pp_28_16, s323, c323);
    logic s324 ,c324; 
    fa fa324 (pp_29_14, pp_30_12, pp_31_10, s324, c324);
    logic s325 ,c325; 
    fa fa325 (c59, c60, s61, s325, c325);
    logic s326 ,c326; 
    fa fa326 (pp_7_59, pp_8_57, pp_9_55, s326, c326);
    logic s327 ,c327; 
    fa fa327 (pp_10_53, pp_11_51, pp_12_49, s327, c327);
    logic s328 ,c328; 
    fa fa328 (pp_13_47, pp_14_45, pp_15_43, s328, c328);
    logic s329 ,c329; 
    fa fa329 (pp_16_41, pp_17_39, pp_18_37, s329, c329);
    logic s330 ,c330; 
    fa fa330 (pp_19_35, pp_20_33, pp_21_31, s330, c330);
    logic s331 ,c331; 
    fa fa331 (pp_22_29, pp_23_27, pp_24_25, s331, c331);
    logic s332 ,c332; 
    fa fa332 (pp_25_23, pp_26_21, pp_27_19, s332, c332);
    logic s333 ,c333; 
    fa fa333 (pp_28_17, pp_29_15, pp_30_13, s333, c333);
    logic s334 ,c334; 
    fa fa334 (pp_31_11, c61, c62, s334, c334);
    logic s335 ,c335; 
    fa fa335 (pp_6_62, pp_7_60, pp_8_58, s335, c335);
    logic s336 ,c336; 
    fa fa336 (pp_9_56, pp_10_54, pp_11_52, s336, c336);
    logic s337 ,c337; 
    fa fa337 (pp_12_50, pp_13_48, pp_14_46, s337, c337);
    logic s338 ,c338; 
    fa fa338 (pp_15_44, pp_16_42, pp_17_40, s338, c338);
    logic s339 ,c339; 
    fa fa339 (pp_18_38, pp_19_36, pp_20_34, s339, c339);
    logic s340 ,c340; 
    fa fa340 (pp_21_32, pp_22_30, pp_23_28, s340, c340);
    logic s341 ,c341; 
    fa fa341 (pp_24_26, pp_25_24, pp_26_22, s341, c341);
    logic s342 ,c342; 
    fa fa342 (pp_27_20, pp_28_18, pp_29_16, s342, c342);
    logic s343 ,c343; 
    fa fa343 (pp_30_14, pp_31_12, c63, s343, c343);
    logic s344 ,c344; 
    fa fa344 (pp_5_65, pp_6_63, pp_7_61, s344, c344);
    logic s345 ,c345; 
    fa fa345 (pp_8_59, pp_9_57, pp_10_55, s345, c345);
    logic s346 ,c346; 
    fa fa346 (pp_11_53, pp_12_51, pp_13_49, s346, c346);
    logic s347 ,c347; 
    fa fa347 (pp_14_47, pp_15_45, pp_16_43, s347, c347);
    logic s348 ,c348; 
    fa fa348 (pp_17_41, pp_18_39, pp_19_37, s348, c348);
    logic s349 ,c349; 
    fa fa349 (pp_20_35, pp_21_33, pp_22_31, s349, c349);
    logic s350 ,c350; 
    fa fa350 (pp_23_29, pp_24_27, pp_25_25, s350, c350);
    logic s351 ,c351; 
    fa fa351 (pp_26_23, pp_27_21, pp_28_19, s351, c351);
    logic s352 ,c352; 
    fa fa352 (pp_29_17, pp_30_15, pp_31_13, s352, c352);
    logic s353 ,c353; 
    fa fa353 (const1, pp_6_64, pp_7_62, s353, c353);
    logic s354 ,c354; 
    fa fa354 (pp_8_60, pp_9_58, pp_10_56, s354, c354);
    logic s355 ,c355; 
    fa fa355 (pp_11_54, pp_12_52, pp_13_50, s355, c355);
    logic s356 ,c356; 
    fa fa356 (pp_14_48, pp_15_46, pp_16_44, s356, c356);
    logic s357 ,c357; 
    fa fa357 (pp_17_42, pp_18_40, pp_19_38, s357, c357);
    logic s358 ,c358; 
    fa fa358 (pp_20_36, pp_21_34, pp_22_32, s358, c358);
    logic s359 ,c359; 
    fa fa359 (pp_23_30, pp_24_28, pp_25_26, s359, c359);
    logic s360 ,c360; 
    fa fa360 (pp_26_24, pp_27_22, pp_28_20, s360, c360);
    logic s361 ,c361;
    ha ha361 (pp_29_18, pp_30_16, s361, c361);
    logic s362 ,c362; 
    fa fa362 (pp_6_65, pp_7_63, pp_8_61, s362, c362);
    logic s363 ,c363; 
    fa fa363 (pp_9_59, pp_10_57, pp_11_55, s363, c363);
    logic s364 ,c364; 
    fa fa364 (pp_12_53, pp_13_51, pp_14_49, s364, c364);
    logic s365 ,c365; 
    fa fa365 (pp_15_47, pp_16_45, pp_17_43, s365, c365);
    logic s366 ,c366; 
    fa fa366 (pp_18_41, pp_19_39, pp_20_37, s366, c366);
    logic s367 ,c367; 
    fa fa367 (pp_21_35, pp_22_33, pp_23_31, s367, c367);
    logic s368 ,c368; 
    fa fa368 (pp_24_29, pp_25_27, pp_26_25, s368, c368);
    logic s369 ,c369; 
    fa fa369 (pp_27_23, pp_28_21, pp_29_19, s369, c369);
    logic s370 ,c370; 
    fa fa370 (const1, pp_7_64, pp_8_62, s370, c370);
    logic s371 ,c371; 
    fa fa371 (pp_9_60, pp_10_58, pp_11_56, s371, c371);
    logic s372 ,c372; 
    fa fa372 (pp_12_54, pp_13_52, pp_14_50, s372, c372);
    logic s373 ,c373; 
    fa fa373 (pp_15_48, pp_16_46, pp_17_44, s373, c373);
    logic s374 ,c374; 
    fa fa374 (pp_18_42, pp_19_40, pp_20_38, s374, c374);
    logic s375 ,c375; 
    fa fa375 (pp_21_36, pp_22_34, pp_23_32, s375, c375);
    logic s376 ,c376; 
    fa fa376 (pp_24_30, pp_25_28, pp_26_26, s376, c376);
    logic s377 ,c377;
    ha ha377 (pp_27_24, pp_28_22, s377, c377);
    logic s378 ,c378; 
    fa fa378 (pp_7_65, pp_8_63, pp_9_61, s378, c378);
    logic s379 ,c379; 
    fa fa379 (pp_10_59, pp_11_57, pp_12_55, s379, c379);
    logic s380 ,c380; 
    fa fa380 (pp_13_53, pp_14_51, pp_15_49, s380, c380);
    logic s381 ,c381; 
    fa fa381 (pp_16_47, pp_17_45, pp_18_43, s381, c381);
    logic s382 ,c382; 
    fa fa382 (pp_19_41, pp_20_39, pp_21_37, s382, c382);
    logic s383 ,c383; 
    fa fa383 (pp_22_35, pp_23_33, pp_24_31, s383, c383);
    logic s384 ,c384; 
    fa fa384 (pp_25_29, pp_26_27, pp_27_25, s384, c384);
    logic s385 ,c385; 
    fa fa385 (const1, pp_8_64, pp_9_62, s385, c385);
    logic s386 ,c386; 
    fa fa386 (pp_10_60, pp_11_58, pp_12_56, s386, c386);
    logic s387 ,c387; 
    fa fa387 (pp_13_54, pp_14_52, pp_15_50, s387, c387);
    logic s388 ,c388; 
    fa fa388 (pp_16_48, pp_17_46, pp_18_44, s388, c388);
    logic s389 ,c389; 
    fa fa389 (pp_19_42, pp_20_40, pp_21_38, s389, c389);
    logic s390 ,c390; 
    fa fa390 (pp_22_36, pp_23_34, pp_24_32, s390, c390);
    logic s391 ,c391;
    ha ha391 (pp_25_30, pp_26_28, s391, c391);
    logic s392 ,c392; 
    fa fa392 (pp_8_65, pp_9_63, pp_10_61, s392, c392);
    logic s393 ,c393; 
    fa fa393 (pp_11_59, pp_12_57, pp_13_55, s393, c393);
    logic s394 ,c394; 
    fa fa394 (pp_14_53, pp_15_51, pp_16_49, s394, c394);
    logic s395 ,c395; 
    fa fa395 (pp_17_47, pp_18_45, pp_19_43, s395, c395);
    logic s396 ,c396; 
    fa fa396 (pp_20_41, pp_21_39, pp_22_37, s396, c396);
    logic s397 ,c397; 
    fa fa397 (pp_23_35, pp_24_33, pp_25_31, s397, c397);
    logic s398 ,c398; 
    fa fa398 (const1, pp_9_64, pp_10_62, s398, c398);
    logic s399 ,c399; 
    fa fa399 (pp_11_60, pp_12_58, pp_13_56, s399, c399);
    logic s400 ,c400; 
    fa fa400 (pp_14_54, pp_15_52, pp_16_50, s400, c400);
    logic s401 ,c401; 
    fa fa401 (pp_17_48, pp_18_46, pp_19_44, s401, c401);
    logic s402 ,c402; 
    fa fa402 (pp_20_42, pp_21_40, pp_22_38, s402, c402);
    logic s403 ,c403;
    ha ha403 (pp_23_36, pp_24_34, s403, c403);
    logic s404 ,c404; 
    fa fa404 (pp_9_65, pp_10_63, pp_11_61, s404, c404);
    logic s405 ,c405; 
    fa fa405 (pp_12_59, pp_13_57, pp_14_55, s405, c405);
    logic s406 ,c406; 
    fa fa406 (pp_15_53, pp_16_51, pp_17_49, s406, c406);
    logic s407 ,c407; 
    fa fa407 (pp_18_47, pp_19_45, pp_20_43, s407, c407);
    logic s408 ,c408; 
    fa fa408 (pp_21_41, pp_22_39, pp_23_37, s408, c408);
    logic s409 ,c409; 
    fa fa409 (const1, pp_10_64, pp_11_62, s409, c409);
    logic s410 ,c410; 
    fa fa410 (pp_12_60, pp_13_58, pp_14_56, s410, c410);
    logic s411 ,c411; 
    fa fa411 (pp_15_54, pp_16_52, pp_17_50, s411, c411);
    logic s412 ,c412; 
    fa fa412 (pp_18_48, pp_19_46, pp_20_44, s412, c412);
    logic s413 ,c413;
    ha ha413 (pp_21_42, pp_22_40, s413, c413);
    logic s414 ,c414; 
    fa fa414 (pp_10_65, pp_11_63, pp_12_61, s414, c414);
    logic s415 ,c415; 
    fa fa415 (pp_13_59, pp_14_57, pp_15_55, s415, c415);
    logic s416 ,c416; 
    fa fa416 (pp_16_53, pp_17_51, pp_18_49, s416, c416);
    logic s417 ,c417; 
    fa fa417 (pp_19_47, pp_20_45, pp_21_43, s417, c417);
    logic s418 ,c418; 
    fa fa418 (const1, pp_11_64, pp_12_62, s418, c418);
    logic s419 ,c419; 
    fa fa419 (pp_13_60, pp_14_58, pp_15_56, s419, c419);
    logic s420 ,c420; 
    fa fa420 (pp_16_54, pp_17_52, pp_18_50, s420, c420);
    logic s421 ,c421;
    ha ha421 (pp_19_48, pp_20_46, s421, c421);
    logic s422 ,c422; 
    fa fa422 (pp_11_65, pp_12_63, pp_13_61, s422, c422);
    logic s423 ,c423; 
    fa fa423 (pp_14_59, pp_15_57, pp_16_55, s423, c423);
    logic s424 ,c424; 
    fa fa424 (pp_17_53, pp_18_51, pp_19_49, s424, c424);
    logic s425 ,c425; 
    fa fa425 (const1, pp_12_64, pp_13_62, s425, c425);
    logic s426 ,c426; 
    fa fa426 (pp_14_60, pp_15_58, pp_16_56, s426, c426);
    logic s427 ,c427;
    ha ha427 (pp_17_54, pp_18_52, s427, c427);
    logic s428 ,c428; 
    fa fa428 (pp_12_65, pp_13_63, pp_14_61, s428, c428);
    logic s429 ,c429; 
    fa fa429 (pp_15_59, pp_16_57, pp_17_55, s429, c429);
    logic s430 ,c430; 
    fa fa430 (const1, pp_13_64, pp_14_62, s430, c430);
    logic s431 ,c431;
    ha ha431 (pp_15_60, pp_16_58, s431, c431);
    logic s432 ,c432; 
    fa fa432 (pp_13_65, pp_14_63, pp_15_61, s432, c432);
    logic s433 ,c433;
    ha ha433 (const1, pp_14_64, s433, c433);
    logic s434 ,c434;
    ha ha434 (pp_0_24, pp_1_22, s434, c434);
    logic s435 ,c435;
    ha ha435 (pp_0_25, pp_1_23, s435, c435);
    logic s436 ,c436; 
    fa fa436 (pp_0_26, pp_1_24, pp_2_22, s436, c436);
    logic s437 ,c437;
    ha ha437 (pp_3_20, pp_4_18, s437, c437);
    logic s438 ,c438; 
    fa fa438 (pp_0_27, pp_1_25, pp_2_23, s438, c438);
    logic s439 ,c439;
    ha ha439 (pp_3_21, pp_4_19, s439, c439);
    logic s440 ,c440; 
    fa fa440 (pp_0_28, pp_1_26, pp_2_24, s440, c440);
    logic s441 ,c441; 
    fa fa441 (pp_3_22, pp_4_20, pp_5_18, s441, c441);
    logic s442 ,c442;
    ha ha442 (pp_6_16, pp_7_14, s442, c442);
    logic s443 ,c443; 
    fa fa443 (pp_0_29, pp_1_27, pp_2_25, s443, c443);
    logic s444 ,c444; 
    fa fa444 (pp_3_23, pp_4_21, pp_5_19, s444, c444);
    logic s445 ,c445;
    ha ha445 (pp_6_17, pp_7_15, s445, c445);
    logic s446 ,c446; 
    fa fa446 (pp_0_30, pp_1_28, pp_2_26, s446, c446);
    logic s447 ,c447; 
    fa fa447 (pp_3_24, pp_4_22, pp_5_20, s447, c447);
    logic s448 ,c448; 
    fa fa448 (pp_6_18, pp_7_16, pp_8_14, s448, c448);
    logic s449 ,c449;
    ha ha449 (pp_9_12, pp_10_10, s449, c449);
    logic s450 ,c450; 
    fa fa450 (pp_0_31, pp_1_29, pp_2_27, s450, c450);
    logic s451 ,c451; 
    fa fa451 (pp_3_25, pp_4_23, pp_5_21, s451, c451);
    logic s452 ,c452; 
    fa fa452 (pp_6_19, pp_7_17, pp_8_15, s452, c452);
    logic s453 ,c453;
    ha ha453 (pp_9_13, pp_10_11, s453, c453);
    logic s454 ,c454; 
    fa fa454 (pp_0_32, pp_1_30, pp_2_28, s454, c454);
    logic s455 ,c455; 
    fa fa455 (pp_3_26, pp_4_24, pp_5_22, s455, c455);
    logic s456 ,c456; 
    fa fa456 (pp_6_20, pp_7_18, pp_8_16, s456, c456);
    logic s457 ,c457; 
    fa fa457 (pp_9_14, pp_10_12, pp_11_10, s457, c457);
    logic s458 ,c458;
    ha ha458 (pp_12_8, pp_13_6, s458, c458);
    logic s459 ,c459; 
    fa fa459 (pp_0_33, pp_1_31, pp_2_29, s459, c459);
    logic s460 ,c460; 
    fa fa460 (pp_3_27, pp_4_25, pp_5_23, s460, c460);
    logic s461 ,c461; 
    fa fa461 (pp_6_21, pp_7_19, pp_8_17, s461, c461);
    logic s462 ,c462; 
    fa fa462 (pp_9_15, pp_10_13, pp_11_11, s462, c462);
    logic s463 ,c463;
    ha ha463 (pp_12_9, pp_13_7, s463, c463);
    logic s464 ,c464; 
    fa fa464 (pp_0_34, pp_1_32, pp_2_30, s464, c464);
    logic s465 ,c465; 
    fa fa465 (pp_3_28, pp_4_26, pp_5_24, s465, c465);
    logic s466 ,c466; 
    fa fa466 (pp_6_22, pp_7_20, pp_8_18, s466, c466);
    logic s467 ,c467; 
    fa fa467 (pp_9_16, pp_10_14, pp_11_12, s467, c467);
    logic s468 ,c468; 
    fa fa468 (pp_12_10, pp_13_8, pp_14_6, s468, c468);
    logic s469 ,c469;
    ha ha469 (pp_15_4, pp_16_2, s469, c469);
    logic s470 ,c470; 
    fa fa470 (pp_0_35, pp_1_33, pp_2_31, s470, c470);
    logic s471 ,c471; 
    fa fa471 (pp_3_29, pp_4_27, pp_5_25, s471, c471);
    logic s472 ,c472; 
    fa fa472 (pp_6_23, pp_7_21, pp_8_19, s472, c472);
    logic s473 ,c473; 
    fa fa473 (pp_9_17, pp_10_15, pp_11_13, s473, c473);
    logic s474 ,c474; 
    fa fa474 (pp_12_11, pp_13_9, pp_14_7, s474, c474);
    logic s475 ,c475;
    ha ha475 (pp_15_5, pp_16_3, s475, c475);
    logic s476 ,c476; 
    fa fa476 (pp_2_32, pp_3_30, pp_4_28, s476, c476);
    logic s477 ,c477; 
    fa fa477 (pp_5_26, pp_6_24, pp_7_22, s477, c477);
    logic s478 ,c478; 
    fa fa478 (pp_8_20, pp_9_18, pp_10_16, s478, c478);
    logic s479 ,c479; 
    fa fa479 (pp_11_14, pp_12_12, pp_13_10, s479, c479);
    logic s480 ,c480; 
    fa fa480 (pp_14_8, pp_15_6, pp_16_4, s480, c480);
    logic s481 ,c481; 
    fa fa481 (pp_17_2, pp_18_0, tcomp18, s481, c481);
    logic s482 ,c482; 
    fa fa482 (pp_2_33, pp_3_31, pp_4_29, s482, c482);
    logic s483 ,c483; 
    fa fa483 (pp_5_27, pp_6_25, pp_7_23, s483, c483);
    logic s484 ,c484; 
    fa fa484 (pp_8_21, pp_9_19, pp_10_17, s484, c484);
    logic s485 ,c485; 
    fa fa485 (pp_11_15, pp_12_13, pp_13_11, s485, c485);
    logic s486 ,c486; 
    fa fa486 (pp_14_9, pp_15_7, pp_16_5, s486, c486);
    logic s487 ,c487; 
    fa fa487 (pp_17_3, pp_18_1, c65, s487, c487);
    logic s488 ,c488; 
    fa fa488 (pp_5_28, pp_6_26, pp_7_24, s488, c488);
    logic s489 ,c489; 
    fa fa489 (pp_8_22, pp_9_20, pp_10_18, s489, c489);
    logic s490 ,c490; 
    fa fa490 (pp_11_16, pp_12_14, pp_13_12, s490, c490);
    logic s491 ,c491; 
    fa fa491 (pp_14_10, pp_15_8, pp_16_6, s491, c491);
    logic s492 ,c492; 
    fa fa492 (pp_17_4, pp_18_2, pp_19_0, s492, c492);
    logic s493 ,c493; 
    fa fa493 (tcomp19, c66, s67, s493, c493);
    logic s494 ,c494; 
    fa fa494 (pp_5_29, pp_6_27, pp_7_25, s494, c494);
    logic s495 ,c495; 
    fa fa495 (pp_8_23, pp_9_21, pp_10_19, s495, c495);
    logic s496 ,c496; 
    fa fa496 (pp_11_17, pp_12_15, pp_13_13, s496, c496);
    logic s497 ,c497; 
    fa fa497 (pp_14_11, pp_15_9, pp_16_7, s497, c497);
    logic s498 ,c498; 
    fa fa498 (pp_17_5, pp_18_3, pp_19_1, s498, c498);
    logic s499 ,c499; 
    fa fa499 (c67, c68, s69, s499, c499);
    logic s500 ,c500; 
    fa fa500 (pp_8_24, pp_9_22, pp_10_20, s500, c500);
    logic s501 ,c501; 
    fa fa501 (pp_11_18, pp_12_16, pp_13_14, s501, c501);
    logic s502 ,c502; 
    fa fa502 (pp_14_12, pp_15_10, pp_16_8, s502, c502);
    logic s503 ,c503; 
    fa fa503 (pp_17_6, pp_18_4, pp_19_2, s503, c503);
    logic s504 ,c504; 
    fa fa504 (pp_20_0, tcomp20, c69, s504, c504);
    logic s505 ,c505; 
    fa fa505 (c70, s71, s72, s505, c505);
    logic s506 ,c506; 
    fa fa506 (pp_8_25, pp_9_23, pp_10_21, s506, c506);
    logic s507 ,c507; 
    fa fa507 (pp_11_19, pp_12_17, pp_13_15, s507, c507);
    logic s508 ,c508; 
    fa fa508 (pp_14_13, pp_15_11, pp_16_9, s508, c508);
    logic s509 ,c509; 
    fa fa509 (pp_17_7, pp_18_5, pp_19_3, s509, c509);
    logic s510 ,c510; 
    fa fa510 (pp_20_1, c71, c72, s510, c510);
    logic s511 ,c511; 
    fa fa511 (c73, s74, s75, s511, c511);
    logic s512 ,c512; 
    fa fa512 (pp_11_20, pp_12_18, pp_13_16, s512, c512);
    logic s513 ,c513; 
    fa fa513 (pp_14_14, pp_15_12, pp_16_10, s513, c513);
    logic s514 ,c514; 
    fa fa514 (pp_17_8, pp_18_6, pp_19_4, s514, c514);
    logic s515 ,c515; 
    fa fa515 (pp_20_2, pp_21_0, tcomp21, s515, c515);
    logic s516 ,c516; 
    fa fa516 (c74, c75, c76, s516, c516);
    logic s517 ,c517; 
    fa fa517 (s77, s78, s79, s517, c517);
    logic s518 ,c518; 
    fa fa518 (pp_11_21, pp_12_19, pp_13_17, s518, c518);
    logic s519 ,c519; 
    fa fa519 (pp_14_15, pp_15_13, pp_16_11, s519, c519);
    logic s520 ,c520; 
    fa fa520 (pp_17_9, pp_18_7, pp_19_5, s520, c520);
    logic s521 ,c521; 
    fa fa521 (pp_20_3, pp_21_1, c77, s521, c521);
    logic s522 ,c522; 
    fa fa522 (c78, c79, c80, s522, c522);
    logic s523 ,c523; 
    fa fa523 (s81, s82, s83, s523, c523);
    logic s524 ,c524; 
    fa fa524 (pp_14_16, pp_15_14, pp_16_12, s524, c524);
    logic s525 ,c525; 
    fa fa525 (pp_17_10, pp_18_8, pp_19_6, s525, c525);
    logic s526 ,c526; 
    fa fa526 (pp_20_4, pp_21_2, pp_22_0, s526, c526);
    logic s527 ,c527; 
    fa fa527 (tcomp22, c81, c82, s527, c527);
    logic s528 ,c528; 
    fa fa528 (c83, c84, s85, s528, c528);
    logic s529 ,c529; 
    fa fa529 (s86, s87, s88, s529, c529);
    logic s530 ,c530; 
    fa fa530 (pp_14_17, pp_15_15, pp_16_13, s530, c530);
    logic s531 ,c531; 
    fa fa531 (pp_17_11, pp_18_9, pp_19_7, s531, c531);
    logic s532 ,c532; 
    fa fa532 (pp_20_5, pp_21_3, pp_22_1, s532, c532);
    logic s533 ,c533; 
    fa fa533 (c85, c86, c87, s533, c533);
    logic s534 ,c534; 
    fa fa534 (c88, c89, s90, s534, c534);
    logic s535 ,c535; 
    fa fa535 (s91, s92, s93, s535, c535);
    logic s536 ,c536; 
    fa fa536 (pp_17_12, pp_18_10, pp_19_8, s536, c536);
    logic s537 ,c537; 
    fa fa537 (pp_20_6, pp_21_4, pp_22_2, s537, c537);
    logic s538 ,c538; 
    fa fa538 (pp_23_0, tcomp23, c90, s538, c538);
    logic s539 ,c539; 
    fa fa539 (c91, c92, c93, s539, c539);
    logic s540 ,c540; 
    fa fa540 (c94, s95, s96, s540, c540);
    logic s541 ,c541; 
    fa fa541 (s97, s98, s99, s541, c541);
    logic s542 ,c542; 
    fa fa542 (pp_17_13, pp_18_11, pp_19_9, s542, c542);
    logic s543 ,c543; 
    fa fa543 (pp_20_7, pp_21_5, pp_22_3, s543, c543);
    logic s544 ,c544; 
    fa fa544 (pp_23_1, c95, c96, s544, c544);
    logic s545 ,c545; 
    fa fa545 (c97, c98, c99, s545, c545);
    logic s546 ,c546; 
    fa fa546 (c100, s101, s102, s546, c546);
    logic s547 ,c547; 
    fa fa547 (s103, s104, s105, s547, c547);
    logic s548 ,c548; 
    fa fa548 (pp_20_8, pp_21_6, pp_22_4, s548, c548);
    logic s549 ,c549; 
    fa fa549 (pp_23_2, pp_24_0, tcomp24, s549, c549);
    logic s550 ,c550; 
    fa fa550 (c101, c102, c103, s550, c550);
    logic s551 ,c551; 
    fa fa551 (c104, c105, c106, s551, c551);
    logic s552 ,c552; 
    fa fa552 (s107, s108, s109, s552, c552);
    logic s553 ,c553; 
    fa fa553 (s110, s111, s112, s553, c553);
    logic s554 ,c554; 
    fa fa554 (pp_20_9, pp_21_7, pp_22_5, s554, c554);
    logic s555 ,c555; 
    fa fa555 (pp_23_3, pp_24_1, c107, s555, c555);
    logic s556 ,c556; 
    fa fa556 (c108, c109, c110, s556, c556);
    logic s557 ,c557; 
    fa fa557 (c111, c112, c113, s557, c557);
    logic s558 ,c558; 
    fa fa558 (s114, s115, s116, s558, c558);
    logic s559 ,c559; 
    fa fa559 (s117, s118, s119, s559, c559);
    logic s560 ,c560; 
    fa fa560 (pp_23_4, pp_24_2, pp_25_0, s560, c560);
    logic s561 ,c561; 
    fa fa561 (tcomp25, c114, c115, s561, c561);
    logic s562 ,c562; 
    fa fa562 (c116, c117, c118, s562, c562);
    logic s563 ,c563; 
    fa fa563 (c119, c120, s121, s563, c563);
    logic s564 ,c564; 
    fa fa564 (s122, s123, s124, s564, c564);
    logic s565 ,c565; 
    fa fa565 (s125, s126, s127, s565, c565);
    logic s566 ,c566; 
    fa fa566 (pp_23_5, pp_24_3, pp_25_1, s566, c566);
    logic s567 ,c567; 
    fa fa567 (c121, c122, c123, s567, c567);
    logic s568 ,c568; 
    fa fa568 (c124, c125, c126, s568, c568);
    logic s569 ,c569; 
    fa fa569 (c127, c128, s129, s569, c569);
    logic s570 ,c570; 
    fa fa570 (s130, s131, s132, s570, c570);
    logic s571 ,c571; 
    fa fa571 (s133, s134, s135, s571, c571);
    logic s572 ,c572; 
    fa fa572 (pp_26_0, tcomp26, c129, s572, c572);
    logic s573 ,c573; 
    fa fa573 (c130, c131, c132, s573, c573);
    logic s574 ,c574; 
    fa fa574 (c133, c134, c135, s574, c574);
    logic s575 ,c575; 
    fa fa575 (c136, s137, s138, s575, c575);
    logic s576 ,c576; 
    fa fa576 (s139, s140, s141, s576, c576);
    logic s577 ,c577; 
    fa fa577 (s142, s143, s144, s577, c577);
    logic s578 ,c578; 
    fa fa578 (pp_26_1, c137, c138, s578, c578);
    logic s579 ,c579; 
    fa fa579 (c139, c140, c141, s579, c579);
    logic s580 ,c580; 
    fa fa580 (c142, c143, c144, s580, c580);
    logic s581 ,c581; 
    fa fa581 (c145, s146, s147, s581, c581);
    logic s582 ,c582; 
    fa fa582 (s148, s149, s150, s582, c582);
    logic s583 ,c583; 
    fa fa583 (s151, s152, s153, s583, c583);
    logic s584 ,c584; 
    fa fa584 (s0, c146, c147, s584, c584);
    logic s585 ,c585; 
    fa fa585 (c148, c149, c150, s585, c585);
    logic s586 ,c586; 
    fa fa586 (c151, c152, c153, s586, c586);
    logic s587 ,c587; 
    fa fa587 (c154, s155, s156, s587, c587);
    logic s588 ,c588; 
    fa fa588 (s157, s158, s159, s588, c588);
    logic s589 ,c589; 
    fa fa589 (s160, s161, s162, s589, c589);
    logic s590 ,c590; 
    fa fa590 (s1, c155, c156, s590, c590);
    logic s591 ,c591; 
    fa fa591 (c157, c158, c159, s591, c591);
    logic s592 ,c592; 
    fa fa592 (c160, c161, c162, s592, c592);
    logic s593 ,c593; 
    fa fa593 (c163, s164, s165, s593, c593);
    logic s594 ,c594; 
    fa fa594 (s166, s167, s168, s594, c594);
    logic s595 ,c595; 
    fa fa595 (s169, s170, s171, s595, c595);
    logic s596 ,c596; 
    fa fa596 (s3, c164, c165, s596, c596);
    logic s597 ,c597; 
    fa fa597 (c166, c167, c168, s597, c597);
    logic s598 ,c598; 
    fa fa598 (c169, c170, c171, s598, c598);
    logic s599 ,c599; 
    fa fa599 (c172, s173, s174, s599, c599);
    logic s600 ,c600; 
    fa fa600 (s175, s176, s177, s600, c600);
    logic s601 ,c601; 
    fa fa601 (s178, s179, s180, s601, c601);
    logic s602 ,c602; 
    fa fa602 (s5, c173, c174, s602, c602);
    logic s603 ,c603; 
    fa fa603 (c175, c176, c177, s603, c603);
    logic s604 ,c604; 
    fa fa604 (c178, c179, c180, s604, c604);
    logic s605 ,c605; 
    fa fa605 (c181, s182, s183, s605, c605);
    logic s606 ,c606; 
    fa fa606 (s184, s185, s186, s606, c606);
    logic s607 ,c607; 
    fa fa607 (s187, s188, s189, s607, c607);
    logic s608 ,c608; 
    fa fa608 (s8, c182, c183, s608, c608);
    logic s609 ,c609; 
    fa fa609 (c184, c185, c186, s609, c609);
    logic s610 ,c610; 
    fa fa610 (c187, c188, c189, s610, c610);
    logic s611 ,c611; 
    fa fa611 (c190, s191, s192, s611, c611);
    logic s612 ,c612; 
    fa fa612 (s193, s194, s195, s612, c612);
    logic s613 ,c613; 
    fa fa613 (s196, s197, s198, s613, c613);
    logic s614 ,c614; 
    fa fa614 (s11, c191, c192, s614, c614);
    logic s615 ,c615; 
    fa fa615 (c193, c194, c195, s615, c615);
    logic s616 ,c616; 
    fa fa616 (c196, c197, c198, s616, c616);
    logic s617 ,c617; 
    fa fa617 (c199, s200, s201, s617, c617);
    logic s618 ,c618; 
    fa fa618 (s202, s203, s204, s618, c618);
    logic s619 ,c619; 
    fa fa619 (s205, s206, s207, s619, c619);
    logic s620 ,c620; 
    fa fa620 (s15, c200, c201, s620, c620);
    logic s621 ,c621; 
    fa fa621 (c202, c203, c204, s621, c621);
    logic s622 ,c622; 
    fa fa622 (c205, c206, c207, s622, c622);
    logic s623 ,c623; 
    fa fa623 (c208, s209, s210, s623, c623);
    logic s624 ,c624; 
    fa fa624 (s211, s212, s213, s624, c624);
    logic s625 ,c625; 
    fa fa625 (s214, s215, s216, s625, c625);
    logic s626 ,c626; 
    fa fa626 (s19, c209, c210, s626, c626);
    logic s627 ,c627; 
    fa fa627 (c211, c212, c213, s627, c627);
    logic s628 ,c628; 
    fa fa628 (c214, c215, c216, s628, c628);
    logic s629 ,c629; 
    fa fa629 (c217, s218, s219, s629, c629);
    logic s630 ,c630; 
    fa fa630 (s220, s221, s222, s630, c630);
    logic s631 ,c631; 
    fa fa631 (s223, s224, s225, s631, c631);
    logic s632 ,c632; 
    fa fa632 (s24, c218, c219, s632, c632);
    logic s633 ,c633; 
    fa fa633 (c220, c221, c222, s633, c633);
    logic s634 ,c634; 
    fa fa634 (c223, c224, c225, s634, c634);
    logic s635 ,c635; 
    fa fa635 (c226, s227, s228, s635, c635);
    logic s636 ,c636; 
    fa fa636 (s229, s230, s231, s636, c636);
    logic s637 ,c637; 
    fa fa637 (s232, s233, s234, s637, c637);
    logic s638 ,c638; 
    fa fa638 (s29, c227, c228, s638, c638);
    logic s639 ,c639; 
    fa fa639 (c229, c230, c231, s639, c639);
    logic s640 ,c640; 
    fa fa640 (c232, c233, c234, s640, c640);
    logic s641 ,c641; 
    fa fa641 (c235, s236, s237, s641, c641);
    logic s642 ,c642; 
    fa fa642 (s238, s239, s240, s642, c642);
    logic s643 ,c643; 
    fa fa643 (s241, s242, s243, s643, c643);
    logic s644 ,c644; 
    fa fa644 (s34, c236, c237, s644, c644);
    logic s645 ,c645; 
    fa fa645 (c238, c239, c240, s645, c645);
    logic s646 ,c646; 
    fa fa646 (c241, c242, c243, s646, c646);
    logic s647 ,c647; 
    fa fa647 (c244, s245, s246, s647, c647);
    logic s648 ,c648; 
    fa fa648 (s247, s248, s249, s648, c648);
    logic s649 ,c649; 
    fa fa649 (s250, s251, s252, s649, c649);
    logic s650 ,c650; 
    fa fa650 (s39, c245, c246, s650, c650);
    logic s651 ,c651; 
    fa fa651 (c247, c248, c249, s651, c651);
    logic s652 ,c652; 
    fa fa652 (c250, c251, c252, s652, c652);
    logic s653 ,c653; 
    fa fa653 (c253, s254, s255, s653, c653);
    logic s654 ,c654; 
    fa fa654 (s256, s257, s258, s654, c654);
    logic s655 ,c655; 
    fa fa655 (s259, s260, s261, s655, c655);
    logic s656 ,c656; 
    fa fa656 (s44, c254, c255, s656, c656);
    logic s657 ,c657; 
    fa fa657 (c256, c257, c258, s657, c657);
    logic s658 ,c658; 
    fa fa658 (c259, c260, c261, s658, c658);
    logic s659 ,c659; 
    fa fa659 (c262, s263, s264, s659, c659);
    logic s660 ,c660; 
    fa fa660 (s265, s266, s267, s660, c660);
    logic s661 ,c661; 
    fa fa661 (s268, s269, s270, s661, c661);
    logic s662 ,c662; 
    fa fa662 (s48, c263, c264, s662, c662);
    logic s663 ,c663; 
    fa fa663 (c265, c266, c267, s663, c663);
    logic s664 ,c664; 
    fa fa664 (c268, c269, c270, s664, c664);
    logic s665 ,c665; 
    fa fa665 (c271, s272, s273, s665, c665);
    logic s666 ,c666; 
    fa fa666 (s274, s275, s276, s666, c666);
    logic s667 ,c667; 
    fa fa667 (s277, s278, s279, s667, c667);
    logic s668 ,c668; 
    fa fa668 (s52, c272, c273, s668, c668);
    logic s669 ,c669; 
    fa fa669 (c274, c275, c276, s669, c669);
    logic s670 ,c670; 
    fa fa670 (c277, c278, c279, s670, c670);
    logic s671 ,c671; 
    fa fa671 (c280, s281, s282, s671, c671);
    logic s672 ,c672; 
    fa fa672 (s283, s284, s285, s672, c672);
    logic s673 ,c673; 
    fa fa673 (s286, s287, s288, s673, c673);
    logic s674 ,c674; 
    fa fa674 (s55, c281, c282, s674, c674);
    logic s675 ,c675; 
    fa fa675 (c283, c284, c285, s675, c675);
    logic s676 ,c676; 
    fa fa676 (c286, c287, c288, s676, c676);
    logic s677 ,c677; 
    fa fa677 (c289, s290, s291, s677, c677);
    logic s678 ,c678; 
    fa fa678 (s292, s293, s294, s678, c678);
    logic s679 ,c679; 
    fa fa679 (s295, s296, s297, s679, c679);
    logic s680 ,c680; 
    fa fa680 (s58, c290, c291, s680, c680);
    logic s681 ,c681; 
    fa fa681 (c292, c293, c294, s681, c681);
    logic s682 ,c682; 
    fa fa682 (c295, c296, c297, s682, c682);
    logic s683 ,c683; 
    fa fa683 (c298, s299, s300, s683, c683);
    logic s684 ,c684; 
    fa fa684 (s301, s302, s303, s684, c684);
    logic s685 ,c685; 
    fa fa685 (s304, s305, s306, s685, c685);
    logic s686 ,c686; 
    fa fa686 (s60, c299, c300, s686, c686);
    logic s687 ,c687; 
    fa fa687 (c301, c302, c303, s687, c687);
    logic s688 ,c688; 
    fa fa688 (c304, c305, c306, s688, c688);
    logic s689 ,c689; 
    fa fa689 (c307, s308, s309, s689, c689);
    logic s690 ,c690; 
    fa fa690 (s310, s311, s312, s690, c690);
    logic s691 ,c691; 
    fa fa691 (s313, s314, s315, s691, c691);
    logic s692 ,c692; 
    fa fa692 (s62, c308, c309, s692, c692);
    logic s693 ,c693; 
    fa fa693 (c310, c311, c312, s693, c693);
    logic s694 ,c694; 
    fa fa694 (c313, c314, c315, s694, c694);
    logic s695 ,c695; 
    fa fa695 (c316, s317, s318, s695, c695);
    logic s696 ,c696; 
    fa fa696 (s319, s320, s321, s696, c696);
    logic s697 ,c697; 
    fa fa697 (s322, s323, s324, s697, c697);
    logic s698 ,c698; 
    fa fa698 (s63, c317, c318, s698, c698);
    logic s699 ,c699; 
    fa fa699 (c319, c320, c321, s699, c699);
    logic s700 ,c700; 
    fa fa700 (c322, c323, c324, s700, c700);
    logic s701 ,c701; 
    fa fa701 (c325, s326, s327, s701, c701);
    logic s702 ,c702; 
    fa fa702 (s328, s329, s330, s702, c702);
    logic s703 ,c703; 
    fa fa703 (s331, s332, s333, s703, c703);
    logic s704 ,c704; 
    fa fa704 (s64, c326, c327, s704, c704);
    logic s705 ,c705; 
    fa fa705 (c328, c329, c330, s705, c705);
    logic s706 ,c706; 
    fa fa706 (c331, c332, c333, s706, c706);
    logic s707 ,c707; 
    fa fa707 (c334, s335, s336, s707, c707);
    logic s708 ,c708; 
    fa fa708 (s337, s338, s339, s708, c708);
    logic s709 ,c709; 
    fa fa709 (s340, s341, s342, s709, c709);
    logic s710 ,c710; 
    fa fa710 (c64, c335, c336, s710, c710);
    logic s711 ,c711; 
    fa fa711 (c337, c338, c339, s711, c711);
    logic s712 ,c712; 
    fa fa712 (c340, c341, c342, s712, c712);
    logic s713 ,c713; 
    fa fa713 (c343, s344, s345, s713, c713);
    logic s714 ,c714; 
    fa fa714 (s346, s347, s348, s714, c714);
    logic s715 ,c715; 
    fa fa715 (s349, s350, s351, s715, c715);
    logic s716 ,c716; 
    fa fa716 (pp_31_14, c344, c345, s716, c716);
    logic s717 ,c717; 
    fa fa717 (c346, c347, c348, s717, c717);
    logic s718 ,c718; 
    fa fa718 (c349, c350, c351, s718, c718);
    logic s719 ,c719; 
    fa fa719 (c352, s353, s354, s719, c719);
    logic s720 ,c720; 
    fa fa720 (s355, s356, s357, s720, c720);
    logic s721 ,c721; 
    fa fa721 (s358, s359, s360, s721, c721);
    logic s722 ,c722; 
    fa fa722 (pp_30_17, pp_31_15, c353, s722, c722);
    logic s723 ,c723; 
    fa fa723 (c354, c355, c356, s723, c723);
    logic s724 ,c724; 
    fa fa724 (c357, c358, c359, s724, c724);
    logic s725 ,c725; 
    fa fa725 (c360, c361, s362, s725, c725);
    logic s726 ,c726; 
    fa fa726 (s363, s364, s365, s726, c726);
    logic s727 ,c727; 
    fa fa727 (s366, s367, s368, s727, c727);
    logic s728 ,c728; 
    fa fa728 (pp_29_20, pp_30_18, pp_31_16, s728, c728);
    logic s729 ,c729; 
    fa fa729 (c362, c363, c364, s729, c729);
    logic s730 ,c730; 
    fa fa730 (c365, c366, c367, s730, c730);
    logic s731 ,c731; 
    fa fa731 (c368, c369, s370, s731, c731);
    logic s732 ,c732; 
    fa fa732 (s371, s372, s373, s732, c732);
    logic s733 ,c733; 
    fa fa733 (s374, s375, s376, s733, c733);
    logic s734 ,c734; 
    fa fa734 (pp_28_23, pp_29_21, pp_30_19, s734, c734);
    logic s735 ,c735; 
    fa fa735 (pp_31_17, c370, c371, s735, c735);
    logic s736 ,c736; 
    fa fa736 (c372, c373, c374, s736, c736);
    logic s737 ,c737; 
    fa fa737 (c375, c376, c377, s737, c737);
    logic s738 ,c738; 
    fa fa738 (s378, s379, s380, s738, c738);
    logic s739 ,c739; 
    fa fa739 (s381, s382, s383, s739, c739);
    logic s740 ,c740; 
    fa fa740 (pp_27_26, pp_28_24, pp_29_22, s740, c740);
    logic s741 ,c741; 
    fa fa741 (pp_30_20, pp_31_18, c378, s741, c741);
    logic s742 ,c742; 
    fa fa742 (c379, c380, c381, s742, c742);
    logic s743 ,c743; 
    fa fa743 (c382, c383, c384, s743, c743);
    logic s744 ,c744; 
    fa fa744 (s385, s386, s387, s744, c744);
    logic s745 ,c745; 
    fa fa745 (s388, s389, s390, s745, c745);
    logic s746 ,c746; 
    fa fa746 (pp_26_29, pp_27_27, pp_28_25, s746, c746);
    logic s747 ,c747; 
    fa fa747 (pp_29_23, pp_30_21, pp_31_19, s747, c747);
    logic s748 ,c748; 
    fa fa748 (c385, c386, c387, s748, c748);
    logic s749 ,c749; 
    fa fa749 (c388, c389, c390, s749, c749);
    logic s750 ,c750; 
    fa fa750 (c391, s392, s393, s750, c750);
    logic s751 ,c751; 
    fa fa751 (s394, s395, s396, s751, c751);
    logic s752 ,c752; 
    fa fa752 (pp_25_32, pp_26_30, pp_27_28, s752, c752);
    logic s753 ,c753; 
    fa fa753 (pp_28_26, pp_29_24, pp_30_22, s753, c753);
    logic s754 ,c754; 
    fa fa754 (pp_31_20, c392, c393, s754, c754);
    logic s755 ,c755; 
    fa fa755 (c394, c395, c396, s755, c755);
    logic s756 ,c756; 
    fa fa756 (c397, s398, s399, s756, c756);
    logic s757 ,c757; 
    fa fa757 (s400, s401, s402, s757, c757);
    logic s758 ,c758; 
    fa fa758 (pp_24_35, pp_25_33, pp_26_31, s758, c758);
    logic s759 ,c759; 
    fa fa759 (pp_27_29, pp_28_27, pp_29_25, s759, c759);
    logic s760 ,c760; 
    fa fa760 (pp_30_23, pp_31_21, c398, s760, c760);
    logic s761 ,c761; 
    fa fa761 (c399, c400, c401, s761, c761);
    logic s762 ,c762; 
    fa fa762 (c402, c403, s404, s762, c762);
    logic s763 ,c763; 
    fa fa763 (s405, s406, s407, s763, c763);
    logic s764 ,c764; 
    fa fa764 (pp_23_38, pp_24_36, pp_25_34, s764, c764);
    logic s765 ,c765; 
    fa fa765 (pp_26_32, pp_27_30, pp_28_28, s765, c765);
    logic s766 ,c766; 
    fa fa766 (pp_29_26, pp_30_24, pp_31_22, s766, c766);
    logic s767 ,c767; 
    fa fa767 (c404, c405, c406, s767, c767);
    logic s768 ,c768; 
    fa fa768 (c407, c408, s409, s768, c768);
    logic s769 ,c769; 
    fa fa769 (s410, s411, s412, s769, c769);
    logic s770 ,c770; 
    fa fa770 (pp_22_41, pp_23_39, pp_24_37, s770, c770);
    logic s771 ,c771; 
    fa fa771 (pp_25_35, pp_26_33, pp_27_31, s771, c771);
    logic s772 ,c772; 
    fa fa772 (pp_28_29, pp_29_27, pp_30_25, s772, c772);
    logic s773 ,c773; 
    fa fa773 (pp_31_23, c409, c410, s773, c773);
    logic s774 ,c774; 
    fa fa774 (c411, c412, c413, s774, c774);
    logic s775 ,c775; 
    fa fa775 (s414, s415, s416, s775, c775);
    logic s776 ,c776; 
    fa fa776 (pp_21_44, pp_22_42, pp_23_40, s776, c776);
    logic s777 ,c777; 
    fa fa777 (pp_24_38, pp_25_36, pp_26_34, s777, c777);
    logic s778 ,c778; 
    fa fa778 (pp_27_32, pp_28_30, pp_29_28, s778, c778);
    logic s779 ,c779; 
    fa fa779 (pp_30_26, pp_31_24, c414, s779, c779);
    logic s780 ,c780; 
    fa fa780 (c415, c416, c417, s780, c780);
    logic s781 ,c781; 
    fa fa781 (s418, s419, s420, s781, c781);
    logic s782 ,c782; 
    fa fa782 (pp_20_47, pp_21_45, pp_22_43, s782, c782);
    logic s783 ,c783; 
    fa fa783 (pp_23_41, pp_24_39, pp_25_37, s783, c783);
    logic s784 ,c784; 
    fa fa784 (pp_26_35, pp_27_33, pp_28_31, s784, c784);
    logic s785 ,c785; 
    fa fa785 (pp_29_29, pp_30_27, pp_31_25, s785, c785);
    logic s786 ,c786; 
    fa fa786 (c418, c419, c420, s786, c786);
    logic s787 ,c787; 
    fa fa787 (c421, s422, s423, s787, c787);
    logic s788 ,c788; 
    fa fa788 (pp_19_50, pp_20_48, pp_21_46, s788, c788);
    logic s789 ,c789; 
    fa fa789 (pp_22_44, pp_23_42, pp_24_40, s789, c789);
    logic s790 ,c790; 
    fa fa790 (pp_25_38, pp_26_36, pp_27_34, s790, c790);
    logic s791 ,c791; 
    fa fa791 (pp_28_32, pp_29_30, pp_30_28, s791, c791);
    logic s792 ,c792; 
    fa fa792 (pp_31_26, c422, c423, s792, c792);
    logic s793 ,c793; 
    fa fa793 (c424, s425, s426, s793, c793);
    logic s794 ,c794; 
    fa fa794 (pp_18_53, pp_19_51, pp_20_49, s794, c794);
    logic s795 ,c795; 
    fa fa795 (pp_21_47, pp_22_45, pp_23_43, s795, c795);
    logic s796 ,c796; 
    fa fa796 (pp_24_41, pp_25_39, pp_26_37, s796, c796);
    logic s797 ,c797; 
    fa fa797 (pp_27_35, pp_28_33, pp_29_31, s797, c797);
    logic s798 ,c798; 
    fa fa798 (pp_30_29, pp_31_27, c425, s798, c798);
    logic s799 ,c799; 
    fa fa799 (c426, c427, s428, s799, c799);
    logic s800 ,c800; 
    fa fa800 (pp_17_56, pp_18_54, pp_19_52, s800, c800);
    logic s801 ,c801; 
    fa fa801 (pp_20_50, pp_21_48, pp_22_46, s801, c801);
    logic s802 ,c802; 
    fa fa802 (pp_23_44, pp_24_42, pp_25_40, s802, c802);
    logic s803 ,c803; 
    fa fa803 (pp_26_38, pp_27_36, pp_28_34, s803, c803);
    logic s804 ,c804; 
    fa fa804 (pp_29_32, pp_30_30, pp_31_28, s804, c804);
    logic s805 ,c805; 
    fa fa805 (c428, c429, s430, s805, c805);
    logic s806 ,c806; 
    fa fa806 (pp_16_59, pp_17_57, pp_18_55, s806, c806);
    logic s807 ,c807; 
    fa fa807 (pp_19_53, pp_20_51, pp_21_49, s807, c807);
    logic s808 ,c808; 
    fa fa808 (pp_22_47, pp_23_45, pp_24_43, s808, c808);
    logic s809 ,c809; 
    fa fa809 (pp_25_41, pp_26_39, pp_27_37, s809, c809);
    logic s810 ,c810; 
    fa fa810 (pp_28_35, pp_29_33, pp_30_31, s810, c810);
    logic s811 ,c811; 
    fa fa811 (pp_31_29, c430, c431, s811, c811);
    logic s812 ,c812; 
    fa fa812 (pp_15_62, pp_16_60, pp_17_58, s812, c812);
    logic s813 ,c813; 
    fa fa813 (pp_18_56, pp_19_54, pp_20_52, s813, c813);
    logic s814 ,c814; 
    fa fa814 (pp_21_50, pp_22_48, pp_23_46, s814, c814);
    logic s815 ,c815; 
    fa fa815 (pp_24_44, pp_25_42, pp_26_40, s815, c815);
    logic s816 ,c816; 
    fa fa816 (pp_27_38, pp_28_36, pp_29_34, s816, c816);
    logic s817 ,c817; 
    fa fa817 (pp_30_32, pp_31_30, c432, s817, c817);
    logic s818 ,c818; 
    fa fa818 (pp_14_65, pp_15_63, pp_16_61, s818, c818);
    logic s819 ,c819; 
    fa fa819 (pp_17_59, pp_18_57, pp_19_55, s819, c819);
    logic s820 ,c820; 
    fa fa820 (pp_20_53, pp_21_51, pp_22_49, s820, c820);
    logic s821 ,c821; 
    fa fa821 (pp_23_47, pp_24_45, pp_25_43, s821, c821);
    logic s822 ,c822; 
    fa fa822 (pp_26_41, pp_27_39, pp_28_37, s822, c822);
    logic s823 ,c823; 
    fa fa823 (pp_29_35, pp_30_33, pp_31_31, s823, c823);
    logic s824 ,c824; 
    fa fa824 (const1, pp_15_64, pp_16_62, s824, c824);
    logic s825 ,c825; 
    fa fa825 (pp_17_60, pp_18_58, pp_19_56, s825, c825);
    logic s826 ,c826; 
    fa fa826 (pp_20_54, pp_21_52, pp_22_50, s826, c826);
    logic s827 ,c827; 
    fa fa827 (pp_23_48, pp_24_46, pp_25_44, s827, c827);
    logic s828 ,c828; 
    fa fa828 (pp_26_42, pp_27_40, pp_28_38, s828, c828);
    logic s829 ,c829;
    ha ha829 (pp_29_36, pp_30_34, s829, c829);
    logic s830 ,c830; 
    fa fa830 (pp_15_65, pp_16_63, pp_17_61, s830, c830);
    logic s831 ,c831; 
    fa fa831 (pp_18_59, pp_19_57, pp_20_55, s831, c831);
    logic s832 ,c832; 
    fa fa832 (pp_21_53, pp_22_51, pp_23_49, s832, c832);
    logic s833 ,c833; 
    fa fa833 (pp_24_47, pp_25_45, pp_26_43, s833, c833);
    logic s834 ,c834; 
    fa fa834 (pp_27_41, pp_28_39, pp_29_37, s834, c834);
    logic s835 ,c835; 
    fa fa835 (const1, pp_16_64, pp_17_62, s835, c835);
    logic s836 ,c836; 
    fa fa836 (pp_18_60, pp_19_58, pp_20_56, s836, c836);
    logic s837 ,c837; 
    fa fa837 (pp_21_54, pp_22_52, pp_23_50, s837, c837);
    logic s838 ,c838; 
    fa fa838 (pp_24_48, pp_25_46, pp_26_44, s838, c838);
    logic s839 ,c839;
    ha ha839 (pp_27_42, pp_28_40, s839, c839);
    logic s840 ,c840; 
    fa fa840 (pp_16_65, pp_17_63, pp_18_61, s840, c840);
    logic s841 ,c841; 
    fa fa841 (pp_19_59, pp_20_57, pp_21_55, s841, c841);
    logic s842 ,c842; 
    fa fa842 (pp_22_53, pp_23_51, pp_24_49, s842, c842);
    logic s843 ,c843; 
    fa fa843 (pp_25_47, pp_26_45, pp_27_43, s843, c843);
    logic s844 ,c844; 
    fa fa844 (const1, pp_17_64, pp_18_62, s844, c844);
    logic s845 ,c845; 
    fa fa845 (pp_19_60, pp_20_58, pp_21_56, s845, c845);
    logic s846 ,c846; 
    fa fa846 (pp_22_54, pp_23_52, pp_24_50, s846, c846);
    logic s847 ,c847;
    ha ha847 (pp_25_48, pp_26_46, s847, c847);
    logic s848 ,c848; 
    fa fa848 (pp_17_65, pp_18_63, pp_19_61, s848, c848);
    logic s849 ,c849; 
    fa fa849 (pp_20_59, pp_21_57, pp_22_55, s849, c849);
    logic s850 ,c850; 
    fa fa850 (pp_23_53, pp_24_51, pp_25_49, s850, c850);
    logic s851 ,c851; 
    fa fa851 (const1, pp_18_64, pp_19_62, s851, c851);
    logic s852 ,c852; 
    fa fa852 (pp_20_60, pp_21_58, pp_22_56, s852, c852);
    logic s853 ,c853;
    ha ha853 (pp_23_54, pp_24_52, s853, c853);
    logic s854 ,c854; 
    fa fa854 (pp_18_65, pp_19_63, pp_20_61, s854, c854);
    logic s855 ,c855; 
    fa fa855 (pp_21_59, pp_22_57, pp_23_55, s855, c855);
    logic s856 ,c856; 
    fa fa856 (const1, pp_19_64, pp_20_62, s856, c856);
    logic s857 ,c857;
    ha ha857 (pp_21_60, pp_22_58, s857, c857);
    logic s858 ,c858; 
    fa fa858 (pp_19_65, pp_20_63, pp_21_61, s858, c858);
    logic s859 ,c859;
    ha ha859 (const1, pp_20_64, s859, c859);
    logic s860 ,c860;
    ha ha860 (pp_0_16, pp_1_14, s860, c860);
    logic s861 ,c861;
    ha ha861 (pp_0_17, pp_1_15, s861, c861);
    logic s862 ,c862; 
    fa fa862 (pp_0_18, pp_1_16, pp_2_14, s862, c862);
    logic s863 ,c863;
    ha ha863 (pp_3_12, pp_4_10, s863, c863);
    logic s864 ,c864; 
    fa fa864 (pp_0_19, pp_1_17, pp_2_15, s864, c864);
    logic s865 ,c865;
    ha ha865 (pp_3_13, pp_4_11, s865, c865);
    logic s866 ,c866; 
    fa fa866 (pp_0_20, pp_1_18, pp_2_16, s866, c866);
    logic s867 ,c867; 
    fa fa867 (pp_3_14, pp_4_12, pp_5_10, s867, c867);
    logic s868 ,c868;
    ha ha868 (pp_6_8, pp_7_6, s868, c868);
    logic s869 ,c869; 
    fa fa869 (pp_0_21, pp_1_19, pp_2_17, s869, c869);
    logic s870 ,c870; 
    fa fa870 (pp_3_15, pp_4_13, pp_5_11, s870, c870);
    logic s871 ,c871;
    ha ha871 (pp_6_9, pp_7_7, s871, c871);
    logic s872 ,c872; 
    fa fa872 (pp_0_22, pp_1_20, pp_2_18, s872, c872);
    logic s873 ,c873; 
    fa fa873 (pp_3_16, pp_4_14, pp_5_12, s873, c873);
    logic s874 ,c874; 
    fa fa874 (pp_6_10, pp_7_8, pp_8_6, s874, c874);
    logic s875 ,c875;
    ha ha875 (pp_9_4, pp_10_2, s875, c875);
    logic s876 ,c876; 
    fa fa876 (pp_0_23, pp_1_21, pp_2_19, s876, c876);
    logic s877 ,c877; 
    fa fa877 (pp_3_17, pp_4_15, pp_5_13, s877, c877);
    logic s878 ,c878; 
    fa fa878 (pp_6_11, pp_7_9, pp_8_7, s878, c878);
    logic s879 ,c879;
    ha ha879 (pp_9_5, pp_10_3, s879, c879);
    logic s880 ,c880; 
    fa fa880 (pp_2_20, pp_3_18, pp_4_16, s880, c880);
    logic s881 ,c881; 
    fa fa881 (pp_5_14, pp_6_12, pp_7_10, s881, c881);
    logic s882 ,c882; 
    fa fa882 (pp_8_8, pp_9_6, pp_10_4, s882, c882);
    logic s883 ,c883; 
    fa fa883 (pp_11_2, pp_12_0, tcomp12, s883, c883);
    logic s884 ,c884; 
    fa fa884 (pp_2_21, pp_3_19, pp_4_17, s884, c884);
    logic s885 ,c885; 
    fa fa885 (pp_5_15, pp_6_13, pp_7_11, s885, c885);
    logic s886 ,c886; 
    fa fa886 (pp_8_9, pp_9_7, pp_10_5, s886, c886);
    logic s887 ,c887; 
    fa fa887 (pp_11_3, pp_12_1, c434, s887, c887);
    logic s888 ,c888; 
    fa fa888 (pp_5_16, pp_6_14, pp_7_12, s888, c888);
    logic s889 ,c889; 
    fa fa889 (pp_8_10, pp_9_8, pp_10_6, s889, c889);
    logic s890 ,c890; 
    fa fa890 (pp_11_4, pp_12_2, pp_13_0, s890, c890);
    logic s891 ,c891; 
    fa fa891 (tcomp13, c435, s436, s891, c891);
    logic s892 ,c892; 
    fa fa892 (pp_5_17, pp_6_15, pp_7_13, s892, c892);
    logic s893 ,c893; 
    fa fa893 (pp_8_11, pp_9_9, pp_10_7, s893, c893);
    logic s894 ,c894; 
    fa fa894 (pp_11_5, pp_12_3, pp_13_1, s894, c894);
    logic s895 ,c895; 
    fa fa895 (c436, c437, s438, s895, c895);
    logic s896 ,c896; 
    fa fa896 (pp_8_12, pp_9_10, pp_10_8, s896, c896);
    logic s897 ,c897; 
    fa fa897 (pp_11_6, pp_12_4, pp_13_2, s897, c897);
    logic s898 ,c898; 
    fa fa898 (pp_14_0, tcomp14, c438, s898, c898);
    logic s899 ,c899; 
    fa fa899 (c439, s440, s441, s899, c899);
    logic s900 ,c900; 
    fa fa900 (pp_8_13, pp_9_11, pp_10_9, s900, c900);
    logic s901 ,c901; 
    fa fa901 (pp_11_7, pp_12_5, pp_13_3, s901, c901);
    logic s902 ,c902; 
    fa fa902 (pp_14_1, c440, c441, s902, c902);
    logic s903 ,c903; 
    fa fa903 (c442, s443, s444, s903, c903);
    logic s904 ,c904; 
    fa fa904 (pp_11_8, pp_12_6, pp_13_4, s904, c904);
    logic s905 ,c905; 
    fa fa905 (pp_14_2, pp_15_0, tcomp15, s905, c905);
    logic s906 ,c906; 
    fa fa906 (c443, c444, c445, s906, c906);
    logic s907 ,c907; 
    fa fa907 (s446, s447, s448, s907, c907);
    logic s908 ,c908; 
    fa fa908 (pp_11_9, pp_12_7, pp_13_5, s908, c908);
    logic s909 ,c909; 
    fa fa909 (pp_14_3, pp_15_1, c446, s909, c909);
    logic s910 ,c910; 
    fa fa910 (c447, c448, c449, s910, c910);
    logic s911 ,c911; 
    fa fa911 (s450, s451, s452, s911, c911);
    logic s912 ,c912; 
    fa fa912 (pp_14_4, pp_15_2, pp_16_0, s912, c912);
    logic s913 ,c913; 
    fa fa913 (tcomp16, c450, c451, s913, c913);
    logic s914 ,c914; 
    fa fa914 (c452, c453, s454, s914, c914);
    logic s915 ,c915; 
    fa fa915 (s455, s456, s457, s915, c915);
    logic s916 ,c916; 
    fa fa916 (pp_14_5, pp_15_3, pp_16_1, s916, c916);
    logic s917 ,c917; 
    fa fa917 (c454, c455, c456, s917, c917);
    logic s918 ,c918; 
    fa fa918 (c457, c458, s459, s918, c918);
    logic s919 ,c919; 
    fa fa919 (s460, s461, s462, s919, c919);
    logic s920 ,c920; 
    fa fa920 (pp_17_0, tcomp17, c459, s920, c920);
    logic s921 ,c921; 
    fa fa921 (c460, c461, c462, s921, c921);
    logic s922 ,c922; 
    fa fa922 (c463, s464, s465, s922, c922);
    logic s923 ,c923; 
    fa fa923 (s466, s467, s468, s923, c923);
    logic s924 ,c924; 
    fa fa924 (pp_17_1, c464, c465, s924, c924);
    logic s925 ,c925; 
    fa fa925 (c466, c467, c468, s925, c925);
    logic s926 ,c926; 
    fa fa926 (c469, s470, s471, s926, c926);
    logic s927 ,c927; 
    fa fa927 (s472, s473, s474, s927, c927);
    logic s928 ,c928; 
    fa fa928 (s65, c470, c471, s928, c928);
    logic s929 ,c929; 
    fa fa929 (c472, c473, c474, s929, c929);
    logic s930 ,c930; 
    fa fa930 (c475, s476, s477, s930, c930);
    logic s931 ,c931; 
    fa fa931 (s478, s479, s480, s931, c931);
    logic s932 ,c932; 
    fa fa932 (s66, c476, c477, s932, c932);
    logic s933 ,c933; 
    fa fa933 (c478, c479, c480, s933, c933);
    logic s934 ,c934; 
    fa fa934 (c481, s482, s483, s934, c934);
    logic s935 ,c935; 
    fa fa935 (s484, s485, s486, s935, c935);
    logic s936 ,c936; 
    fa fa936 (s68, c482, c483, s936, c936);
    logic s937 ,c937; 
    fa fa937 (c484, c485, c486, s937, c937);
    logic s938 ,c938; 
    fa fa938 (c487, s488, s489, s938, c938);
    logic s939 ,c939; 
    fa fa939 (s490, s491, s492, s939, c939);
    logic s940 ,c940; 
    fa fa940 (s70, c488, c489, s940, c940);
    logic s941 ,c941; 
    fa fa941 (c490, c491, c492, s941, c941);
    logic s942 ,c942; 
    fa fa942 (c493, s494, s495, s942, c942);
    logic s943 ,c943; 
    fa fa943 (s496, s497, s498, s943, c943);
    logic s944 ,c944; 
    fa fa944 (s73, c494, c495, s944, c944);
    logic s945 ,c945; 
    fa fa945 (c496, c497, c498, s945, c945);
    logic s946 ,c946; 
    fa fa946 (c499, s500, s501, s946, c946);
    logic s947 ,c947; 
    fa fa947 (s502, s503, s504, s947, c947);
    logic s948 ,c948; 
    fa fa948 (s76, c500, c501, s948, c948);
    logic s949 ,c949; 
    fa fa949 (c502, c503, c504, s949, c949);
    logic s950 ,c950; 
    fa fa950 (c505, s506, s507, s950, c950);
    logic s951 ,c951; 
    fa fa951 (s508, s509, s510, s951, c951);
    logic s952 ,c952; 
    fa fa952 (s80, c506, c507, s952, c952);
    logic s953 ,c953; 
    fa fa953 (c508, c509, c510, s953, c953);
    logic s954 ,c954; 
    fa fa954 (c511, s512, s513, s954, c954);
    logic s955 ,c955; 
    fa fa955 (s514, s515, s516, s955, c955);
    logic s956 ,c956; 
    fa fa956 (s84, c512, c513, s956, c956);
    logic s957 ,c957; 
    fa fa957 (c514, c515, c516, s957, c957);
    logic s958 ,c958; 
    fa fa958 (c517, s518, s519, s958, c958);
    logic s959 ,c959; 
    fa fa959 (s520, s521, s522, s959, c959);
    logic s960 ,c960; 
    fa fa960 (s89, c518, c519, s960, c960);
    logic s961 ,c961; 
    fa fa961 (c520, c521, c522, s961, c961);
    logic s962 ,c962; 
    fa fa962 (c523, s524, s525, s962, c962);
    logic s963 ,c963; 
    fa fa963 (s526, s527, s528, s963, c963);
    logic s964 ,c964; 
    fa fa964 (s94, c524, c525, s964, c964);
    logic s965 ,c965; 
    fa fa965 (c526, c527, c528, s965, c965);
    logic s966 ,c966; 
    fa fa966 (c529, s530, s531, s966, c966);
    logic s967 ,c967; 
    fa fa967 (s532, s533, s534, s967, c967);
    logic s968 ,c968; 
    fa fa968 (s100, c530, c531, s968, c968);
    logic s969 ,c969; 
    fa fa969 (c532, c533, c534, s969, c969);
    logic s970 ,c970; 
    fa fa970 (c535, s536, s537, s970, c970);
    logic s971 ,c971; 
    fa fa971 (s538, s539, s540, s971, c971);
    logic s972 ,c972; 
    fa fa972 (s106, c536, c537, s972, c972);
    logic s973 ,c973; 
    fa fa973 (c538, c539, c540, s973, c973);
    logic s974 ,c974; 
    fa fa974 (c541, s542, s543, s974, c974);
    logic s975 ,c975; 
    fa fa975 (s544, s545, s546, s975, c975);
    logic s976 ,c976; 
    fa fa976 (s113, c542, c543, s976, c976);
    logic s977 ,c977; 
    fa fa977 (c544, c545, c546, s977, c977);
    logic s978 ,c978; 
    fa fa978 (c547, s548, s549, s978, c978);
    logic s979 ,c979; 
    fa fa979 (s550, s551, s552, s979, c979);
    logic s980 ,c980; 
    fa fa980 (s120, c548, c549, s980, c980);
    logic s981 ,c981; 
    fa fa981 (c550, c551, c552, s981, c981);
    logic s982 ,c982; 
    fa fa982 (c553, s554, s555, s982, c982);
    logic s983 ,c983; 
    fa fa983 (s556, s557, s558, s983, c983);
    logic s984 ,c984; 
    fa fa984 (s128, c554, c555, s984, c984);
    logic s985 ,c985; 
    fa fa985 (c556, c557, c558, s985, c985);
    logic s986 ,c986; 
    fa fa986 (c559, s560, s561, s986, c986);
    logic s987 ,c987; 
    fa fa987 (s562, s563, s564, s987, c987);
    logic s988 ,c988; 
    fa fa988 (s136, c560, c561, s988, c988);
    logic s989 ,c989; 
    fa fa989 (c562, c563, c564, s989, c989);
    logic s990 ,c990; 
    fa fa990 (c565, s566, s567, s990, c990);
    logic s991 ,c991; 
    fa fa991 (s568, s569, s570, s991, c991);
    logic s992 ,c992; 
    fa fa992 (s145, c566, c567, s992, c992);
    logic s993 ,c993; 
    fa fa993 (c568, c569, c570, s993, c993);
    logic s994 ,c994; 
    fa fa994 (c571, s572, s573, s994, c994);
    logic s995 ,c995; 
    fa fa995 (s574, s575, s576, s995, c995);
    logic s996 ,c996; 
    fa fa996 (s154, c572, c573, s996, c996);
    logic s997 ,c997; 
    fa fa997 (c574, c575, c576, s997, c997);
    logic s998 ,c998; 
    fa fa998 (c577, s578, s579, s998, c998);
    logic s999 ,c999; 
    fa fa999 (s580, s581, s582, s999, c999);
    logic s1000 ,c1000; 
    fa fa1000 (s163, c578, c579, s1000, c1000);
    logic s1001 ,c1001; 
    fa fa1001 (c580, c581, c582, s1001, c1001);
    logic s1002 ,c1002; 
    fa fa1002 (c583, s584, s585, s1002, c1002);
    logic s1003 ,c1003; 
    fa fa1003 (s586, s587, s588, s1003, c1003);
    logic s1004 ,c1004; 
    fa fa1004 (s172, c584, c585, s1004, c1004);
    logic s1005 ,c1005; 
    fa fa1005 (c586, c587, c588, s1005, c1005);
    logic s1006 ,c1006; 
    fa fa1006 (c589, s590, s591, s1006, c1006);
    logic s1007 ,c1007; 
    fa fa1007 (s592, s593, s594, s1007, c1007);
    logic s1008 ,c1008; 
    fa fa1008 (s181, c590, c591, s1008, c1008);
    logic s1009 ,c1009; 
    fa fa1009 (c592, c593, c594, s1009, c1009);
    logic s1010 ,c1010; 
    fa fa1010 (c595, s596, s597, s1010, c1010);
    logic s1011 ,c1011; 
    fa fa1011 (s598, s599, s600, s1011, c1011);
    logic s1012 ,c1012; 
    fa fa1012 (s190, c596, c597, s1012, c1012);
    logic s1013 ,c1013; 
    fa fa1013 (c598, c599, c600, s1013, c1013);
    logic s1014 ,c1014; 
    fa fa1014 (c601, s602, s603, s1014, c1014);
    logic s1015 ,c1015; 
    fa fa1015 (s604, s605, s606, s1015, c1015);
    logic s1016 ,c1016; 
    fa fa1016 (s199, c602, c603, s1016, c1016);
    logic s1017 ,c1017; 
    fa fa1017 (c604, c605, c606, s1017, c1017);
    logic s1018 ,c1018; 
    fa fa1018 (c607, s608, s609, s1018, c1018);
    logic s1019 ,c1019; 
    fa fa1019 (s610, s611, s612, s1019, c1019);
    logic s1020 ,c1020; 
    fa fa1020 (s208, c608, c609, s1020, c1020);
    logic s1021 ,c1021; 
    fa fa1021 (c610, c611, c612, s1021, c1021);
    logic s1022 ,c1022; 
    fa fa1022 (c613, s614, s615, s1022, c1022);
    logic s1023 ,c1023; 
    fa fa1023 (s616, s617, s618, s1023, c1023);
    logic s1024 ,c1024; 
    fa fa1024 (s217, c614, c615, s1024, c1024);
    logic s1025 ,c1025; 
    fa fa1025 (c616, c617, c618, s1025, c1025);
    logic s1026 ,c1026; 
    fa fa1026 (c619, s620, s621, s1026, c1026);
    logic s1027 ,c1027; 
    fa fa1027 (s622, s623, s624, s1027, c1027);
    logic s1028 ,c1028; 
    fa fa1028 (s226, c620, c621, s1028, c1028);
    logic s1029 ,c1029; 
    fa fa1029 (c622, c623, c624, s1029, c1029);
    logic s1030 ,c1030; 
    fa fa1030 (c625, s626, s627, s1030, c1030);
    logic s1031 ,c1031; 
    fa fa1031 (s628, s629, s630, s1031, c1031);
    logic s1032 ,c1032; 
    fa fa1032 (s235, c626, c627, s1032, c1032);
    logic s1033 ,c1033; 
    fa fa1033 (c628, c629, c630, s1033, c1033);
    logic s1034 ,c1034; 
    fa fa1034 (c631, s632, s633, s1034, c1034);
    logic s1035 ,c1035; 
    fa fa1035 (s634, s635, s636, s1035, c1035);
    logic s1036 ,c1036; 
    fa fa1036 (s244, c632, c633, s1036, c1036);
    logic s1037 ,c1037; 
    fa fa1037 (c634, c635, c636, s1037, c1037);
    logic s1038 ,c1038; 
    fa fa1038 (c637, s638, s639, s1038, c1038);
    logic s1039 ,c1039; 
    fa fa1039 (s640, s641, s642, s1039, c1039);
    logic s1040 ,c1040; 
    fa fa1040 (s253, c638, c639, s1040, c1040);
    logic s1041 ,c1041; 
    fa fa1041 (c640, c641, c642, s1041, c1041);
    logic s1042 ,c1042; 
    fa fa1042 (c643, s644, s645, s1042, c1042);
    logic s1043 ,c1043; 
    fa fa1043 (s646, s647, s648, s1043, c1043);
    logic s1044 ,c1044; 
    fa fa1044 (s262, c644, c645, s1044, c1044);
    logic s1045 ,c1045; 
    fa fa1045 (c646, c647, c648, s1045, c1045);
    logic s1046 ,c1046; 
    fa fa1046 (c649, s650, s651, s1046, c1046);
    logic s1047 ,c1047; 
    fa fa1047 (s652, s653, s654, s1047, c1047);
    logic s1048 ,c1048; 
    fa fa1048 (s271, c650, c651, s1048, c1048);
    logic s1049 ,c1049; 
    fa fa1049 (c652, c653, c654, s1049, c1049);
    logic s1050 ,c1050; 
    fa fa1050 (c655, s656, s657, s1050, c1050);
    logic s1051 ,c1051; 
    fa fa1051 (s658, s659, s660, s1051, c1051);
    logic s1052 ,c1052; 
    fa fa1052 (s280, c656, c657, s1052, c1052);
    logic s1053 ,c1053; 
    fa fa1053 (c658, c659, c660, s1053, c1053);
    logic s1054 ,c1054; 
    fa fa1054 (c661, s662, s663, s1054, c1054);
    logic s1055 ,c1055; 
    fa fa1055 (s664, s665, s666, s1055, c1055);
    logic s1056 ,c1056; 
    fa fa1056 (s289, c662, c663, s1056, c1056);
    logic s1057 ,c1057; 
    fa fa1057 (c664, c665, c666, s1057, c1057);
    logic s1058 ,c1058; 
    fa fa1058 (c667, s668, s669, s1058, c1058);
    logic s1059 ,c1059; 
    fa fa1059 (s670, s671, s672, s1059, c1059);
    logic s1060 ,c1060; 
    fa fa1060 (s298, c668, c669, s1060, c1060);
    logic s1061 ,c1061; 
    fa fa1061 (c670, c671, c672, s1061, c1061);
    logic s1062 ,c1062; 
    fa fa1062 (c673, s674, s675, s1062, c1062);
    logic s1063 ,c1063; 
    fa fa1063 (s676, s677, s678, s1063, c1063);
    logic s1064 ,c1064; 
    fa fa1064 (s307, c674, c675, s1064, c1064);
    logic s1065 ,c1065; 
    fa fa1065 (c676, c677, c678, s1065, c1065);
    logic s1066 ,c1066; 
    fa fa1066 (c679, s680, s681, s1066, c1066);
    logic s1067 ,c1067; 
    fa fa1067 (s682, s683, s684, s1067, c1067);
    logic s1068 ,c1068; 
    fa fa1068 (s316, c680, c681, s1068, c1068);
    logic s1069 ,c1069; 
    fa fa1069 (c682, c683, c684, s1069, c1069);
    logic s1070 ,c1070; 
    fa fa1070 (c685, s686, s687, s1070, c1070);
    logic s1071 ,c1071; 
    fa fa1071 (s688, s689, s690, s1071, c1071);
    logic s1072 ,c1072; 
    fa fa1072 (s325, c686, c687, s1072, c1072);
    logic s1073 ,c1073; 
    fa fa1073 (c688, c689, c690, s1073, c1073);
    logic s1074 ,c1074; 
    fa fa1074 (c691, s692, s693, s1074, c1074);
    logic s1075 ,c1075; 
    fa fa1075 (s694, s695, s696, s1075, c1075);
    logic s1076 ,c1076; 
    fa fa1076 (s334, c692, c693, s1076, c1076);
    logic s1077 ,c1077; 
    fa fa1077 (c694, c695, c696, s1077, c1077);
    logic s1078 ,c1078; 
    fa fa1078 (c697, s698, s699, s1078, c1078);
    logic s1079 ,c1079; 
    fa fa1079 (s700, s701, s702, s1079, c1079);
    logic s1080 ,c1080; 
    fa fa1080 (s343, c698, c699, s1080, c1080);
    logic s1081 ,c1081; 
    fa fa1081 (c700, c701, c702, s1081, c1081);
    logic s1082 ,c1082; 
    fa fa1082 (c703, s704, s705, s1082, c1082);
    logic s1083 ,c1083; 
    fa fa1083 (s706, s707, s708, s1083, c1083);
    logic s1084 ,c1084; 
    fa fa1084 (s352, c704, c705, s1084, c1084);
    logic s1085 ,c1085; 
    fa fa1085 (c706, c707, c708, s1085, c1085);
    logic s1086 ,c1086; 
    fa fa1086 (c709, s710, s711, s1086, c1086);
    logic s1087 ,c1087; 
    fa fa1087 (s712, s713, s714, s1087, c1087);
    logic s1088 ,c1088; 
    fa fa1088 (s361, c710, c711, s1088, c1088);
    logic s1089 ,c1089; 
    fa fa1089 (c712, c713, c714, s1089, c1089);
    logic s1090 ,c1090; 
    fa fa1090 (c715, s716, s717, s1090, c1090);
    logic s1091 ,c1091; 
    fa fa1091 (s718, s719, s720, s1091, c1091);
    logic s1092 ,c1092; 
    fa fa1092 (s369, c716, c717, s1092, c1092);
    logic s1093 ,c1093; 
    fa fa1093 (c718, c719, c720, s1093, c1093);
    logic s1094 ,c1094; 
    fa fa1094 (c721, s722, s723, s1094, c1094);
    logic s1095 ,c1095; 
    fa fa1095 (s724, s725, s726, s1095, c1095);
    logic s1096 ,c1096; 
    fa fa1096 (s377, c722, c723, s1096, c1096);
    logic s1097 ,c1097; 
    fa fa1097 (c724, c725, c726, s1097, c1097);
    logic s1098 ,c1098; 
    fa fa1098 (c727, s728, s729, s1098, c1098);
    logic s1099 ,c1099; 
    fa fa1099 (s730, s731, s732, s1099, c1099);
    logic s1100 ,c1100; 
    fa fa1100 (s384, c728, c729, s1100, c1100);
    logic s1101 ,c1101; 
    fa fa1101 (c730, c731, c732, s1101, c1101);
    logic s1102 ,c1102; 
    fa fa1102 (c733, s734, s735, s1102, c1102);
    logic s1103 ,c1103; 
    fa fa1103 (s736, s737, s738, s1103, c1103);
    logic s1104 ,c1104; 
    fa fa1104 (s391, c734, c735, s1104, c1104);
    logic s1105 ,c1105; 
    fa fa1105 (c736, c737, c738, s1105, c1105);
    logic s1106 ,c1106; 
    fa fa1106 (c739, s740, s741, s1106, c1106);
    logic s1107 ,c1107; 
    fa fa1107 (s742, s743, s744, s1107, c1107);
    logic s1108 ,c1108; 
    fa fa1108 (s397, c740, c741, s1108, c1108);
    logic s1109 ,c1109; 
    fa fa1109 (c742, c743, c744, s1109, c1109);
    logic s1110 ,c1110; 
    fa fa1110 (c745, s746, s747, s1110, c1110);
    logic s1111 ,c1111; 
    fa fa1111 (s748, s749, s750, s1111, c1111);
    logic s1112 ,c1112; 
    fa fa1112 (s403, c746, c747, s1112, c1112);
    logic s1113 ,c1113; 
    fa fa1113 (c748, c749, c750, s1113, c1113);
    logic s1114 ,c1114; 
    fa fa1114 (c751, s752, s753, s1114, c1114);
    logic s1115 ,c1115; 
    fa fa1115 (s754, s755, s756, s1115, c1115);
    logic s1116 ,c1116; 
    fa fa1116 (s408, c752, c753, s1116, c1116);
    logic s1117 ,c1117; 
    fa fa1117 (c754, c755, c756, s1117, c1117);
    logic s1118 ,c1118; 
    fa fa1118 (c757, s758, s759, s1118, c1118);
    logic s1119 ,c1119; 
    fa fa1119 (s760, s761, s762, s1119, c1119);
    logic s1120 ,c1120; 
    fa fa1120 (s413, c758, c759, s1120, c1120);
    logic s1121 ,c1121; 
    fa fa1121 (c760, c761, c762, s1121, c1121);
    logic s1122 ,c1122; 
    fa fa1122 (c763, s764, s765, s1122, c1122);
    logic s1123 ,c1123; 
    fa fa1123 (s766, s767, s768, s1123, c1123);
    logic s1124 ,c1124; 
    fa fa1124 (s417, c764, c765, s1124, c1124);
    logic s1125 ,c1125; 
    fa fa1125 (c766, c767, c768, s1125, c1125);
    logic s1126 ,c1126; 
    fa fa1126 (c769, s770, s771, s1126, c1126);
    logic s1127 ,c1127; 
    fa fa1127 (s772, s773, s774, s1127, c1127);
    logic s1128 ,c1128; 
    fa fa1128 (s421, c770, c771, s1128, c1128);
    logic s1129 ,c1129; 
    fa fa1129 (c772, c773, c774, s1129, c1129);
    logic s1130 ,c1130; 
    fa fa1130 (c775, s776, s777, s1130, c1130);
    logic s1131 ,c1131; 
    fa fa1131 (s778, s779, s780, s1131, c1131);
    logic s1132 ,c1132; 
    fa fa1132 (s424, c776, c777, s1132, c1132);
    logic s1133 ,c1133; 
    fa fa1133 (c778, c779, c780, s1133, c1133);
    logic s1134 ,c1134; 
    fa fa1134 (c781, s782, s783, s1134, c1134);
    logic s1135 ,c1135; 
    fa fa1135 (s784, s785, s786, s1135, c1135);
    logic s1136 ,c1136; 
    fa fa1136 (s427, c782, c783, s1136, c1136);
    logic s1137 ,c1137; 
    fa fa1137 (c784, c785, c786, s1137, c1137);
    logic s1138 ,c1138; 
    fa fa1138 (c787, s788, s789, s1138, c1138);
    logic s1139 ,c1139; 
    fa fa1139 (s790, s791, s792, s1139, c1139);
    logic s1140 ,c1140; 
    fa fa1140 (s429, c788, c789, s1140, c1140);
    logic s1141 ,c1141; 
    fa fa1141 (c790, c791, c792, s1141, c1141);
    logic s1142 ,c1142; 
    fa fa1142 (c793, s794, s795, s1142, c1142);
    logic s1143 ,c1143; 
    fa fa1143 (s796, s797, s798, s1143, c1143);
    logic s1144 ,c1144; 
    fa fa1144 (s431, c794, c795, s1144, c1144);
    logic s1145 ,c1145; 
    fa fa1145 (c796, c797, c798, s1145, c1145);
    logic s1146 ,c1146; 
    fa fa1146 (c799, s800, s801, s1146, c1146);
    logic s1147 ,c1147; 
    fa fa1147 (s802, s803, s804, s1147, c1147);
    logic s1148 ,c1148; 
    fa fa1148 (s432, c800, c801, s1148, c1148);
    logic s1149 ,c1149; 
    fa fa1149 (c802, c803, c804, s1149, c1149);
    logic s1150 ,c1150; 
    fa fa1150 (c805, s806, s807, s1150, c1150);
    logic s1151 ,c1151; 
    fa fa1151 (s808, s809, s810, s1151, c1151);
    logic s1152 ,c1152; 
    fa fa1152 (s433, c806, c807, s1152, c1152);
    logic s1153 ,c1153; 
    fa fa1153 (c808, c809, c810, s1153, c1153);
    logic s1154 ,c1154; 
    fa fa1154 (c811, s812, s813, s1154, c1154);
    logic s1155 ,c1155; 
    fa fa1155 (s814, s815, s816, s1155, c1155);
    logic s1156 ,c1156; 
    fa fa1156 (c433, c812, c813, s1156, c1156);
    logic s1157 ,c1157; 
    fa fa1157 (c814, c815, c816, s1157, c1157);
    logic s1158 ,c1158; 
    fa fa1158 (c817, s818, s819, s1158, c1158);
    logic s1159 ,c1159; 
    fa fa1159 (s820, s821, s822, s1159, c1159);
    logic s1160 ,c1160; 
    fa fa1160 (pp_31_32, c818, c819, s1160, c1160);
    logic s1161 ,c1161; 
    fa fa1161 (c820, c821, c822, s1161, c1161);
    logic s1162 ,c1162; 
    fa fa1162 (c823, s824, s825, s1162, c1162);
    logic s1163 ,c1163; 
    fa fa1163 (s826, s827, s828, s1163, c1163);
    logic s1164 ,c1164; 
    fa fa1164 (pp_30_35, pp_31_33, c824, s1164, c1164);
    logic s1165 ,c1165; 
    fa fa1165 (c825, c826, c827, s1165, c1165);
    logic s1166 ,c1166; 
    fa fa1166 (c828, c829, s830, s1166, c1166);
    logic s1167 ,c1167; 
    fa fa1167 (s831, s832, s833, s1167, c1167);
    logic s1168 ,c1168; 
    fa fa1168 (pp_29_38, pp_30_36, pp_31_34, s1168, c1168);
    logic s1169 ,c1169; 
    fa fa1169 (c830, c831, c832, s1169, c1169);
    logic s1170 ,c1170; 
    fa fa1170 (c833, c834, s835, s1170, c1170);
    logic s1171 ,c1171; 
    fa fa1171 (s836, s837, s838, s1171, c1171);
    logic s1172 ,c1172; 
    fa fa1172 (pp_28_41, pp_29_39, pp_30_37, s1172, c1172);
    logic s1173 ,c1173; 
    fa fa1173 (pp_31_35, c835, c836, s1173, c1173);
    logic s1174 ,c1174; 
    fa fa1174 (c837, c838, c839, s1174, c1174);
    logic s1175 ,c1175; 
    fa fa1175 (s840, s841, s842, s1175, c1175);
    logic s1176 ,c1176; 
    fa fa1176 (pp_27_44, pp_28_42, pp_29_40, s1176, c1176);
    logic s1177 ,c1177; 
    fa fa1177 (pp_30_38, pp_31_36, c840, s1177, c1177);
    logic s1178 ,c1178; 
    fa fa1178 (c841, c842, c843, s1178, c1178);
    logic s1179 ,c1179; 
    fa fa1179 (s844, s845, s846, s1179, c1179);
    logic s1180 ,c1180; 
    fa fa1180 (pp_26_47, pp_27_45, pp_28_43, s1180, c1180);
    logic s1181 ,c1181; 
    fa fa1181 (pp_29_41, pp_30_39, pp_31_37, s1181, c1181);
    logic s1182 ,c1182; 
    fa fa1182 (c844, c845, c846, s1182, c1182);
    logic s1183 ,c1183; 
    fa fa1183 (c847, s848, s849, s1183, c1183);
    logic s1184 ,c1184; 
    fa fa1184 (pp_25_50, pp_26_48, pp_27_46, s1184, c1184);
    logic s1185 ,c1185; 
    fa fa1185 (pp_28_44, pp_29_42, pp_30_40, s1185, c1185);
    logic s1186 ,c1186; 
    fa fa1186 (pp_31_38, c848, c849, s1186, c1186);
    logic s1187 ,c1187; 
    fa fa1187 (c850, s851, s852, s1187, c1187);
    logic s1188 ,c1188; 
    fa fa1188 (pp_24_53, pp_25_51, pp_26_49, s1188, c1188);
    logic s1189 ,c1189; 
    fa fa1189 (pp_27_47, pp_28_45, pp_29_43, s1189, c1189);
    logic s1190 ,c1190; 
    fa fa1190 (pp_30_41, pp_31_39, c851, s1190, c1190);
    logic s1191 ,c1191; 
    fa fa1191 (c852, c853, s854, s1191, c1191);
    logic s1192 ,c1192; 
    fa fa1192 (pp_23_56, pp_24_54, pp_25_52, s1192, c1192);
    logic s1193 ,c1193; 
    fa fa1193 (pp_26_50, pp_27_48, pp_28_46, s1193, c1193);
    logic s1194 ,c1194; 
    fa fa1194 (pp_29_44, pp_30_42, pp_31_40, s1194, c1194);
    logic s1195 ,c1195; 
    fa fa1195 (c854, c855, s856, s1195, c1195);
    logic s1196 ,c1196; 
    fa fa1196 (pp_22_59, pp_23_57, pp_24_55, s1196, c1196);
    logic s1197 ,c1197; 
    fa fa1197 (pp_25_53, pp_26_51, pp_27_49, s1197, c1197);
    logic s1198 ,c1198; 
    fa fa1198 (pp_28_47, pp_29_45, pp_30_43, s1198, c1198);
    logic s1199 ,c1199; 
    fa fa1199 (pp_31_41, c856, c857, s1199, c1199);
    logic s1200 ,c1200; 
    fa fa1200 (pp_21_62, pp_22_60, pp_23_58, s1200, c1200);
    logic s1201 ,c1201; 
    fa fa1201 (pp_24_56, pp_25_54, pp_26_52, s1201, c1201);
    logic s1202 ,c1202; 
    fa fa1202 (pp_27_50, pp_28_48, pp_29_46, s1202, c1202);
    logic s1203 ,c1203; 
    fa fa1203 (pp_30_44, pp_31_42, c858, s1203, c1203);
    logic s1204 ,c1204; 
    fa fa1204 (pp_20_65, pp_21_63, pp_22_61, s1204, c1204);
    logic s1205 ,c1205; 
    fa fa1205 (pp_23_59, pp_24_57, pp_25_55, s1205, c1205);
    logic s1206 ,c1206; 
    fa fa1206 (pp_26_53, pp_27_51, pp_28_49, s1206, c1206);
    logic s1207 ,c1207; 
    fa fa1207 (pp_29_47, pp_30_45, pp_31_43, s1207, c1207);
    logic s1208 ,c1208; 
    fa fa1208 (const1, pp_21_64, pp_22_62, s1208, c1208);
    logic s1209 ,c1209; 
    fa fa1209 (pp_23_60, pp_24_58, pp_25_56, s1209, c1209);
    logic s1210 ,c1210; 
    fa fa1210 (pp_26_54, pp_27_52, pp_28_50, s1210, c1210);
    logic s1211 ,c1211;
    ha ha1211 (pp_29_48, pp_30_46, s1211, c1211);
    logic s1212 ,c1212; 
    fa fa1212 (pp_21_65, pp_22_63, pp_23_61, s1212, c1212);
    logic s1213 ,c1213; 
    fa fa1213 (pp_24_59, pp_25_57, pp_26_55, s1213, c1213);
    logic s1214 ,c1214; 
    fa fa1214 (pp_27_53, pp_28_51, pp_29_49, s1214, c1214);
    logic s1215 ,c1215; 
    fa fa1215 (const1, pp_22_64, pp_23_62, s1215, c1215);
    logic s1216 ,c1216; 
    fa fa1216 (pp_24_60, pp_25_58, pp_26_56, s1216, c1216);
    logic s1217 ,c1217;
    ha ha1217 (pp_27_54, pp_28_52, s1217, c1217);
    logic s1218 ,c1218; 
    fa fa1218 (pp_22_65, pp_23_63, pp_24_61, s1218, c1218);
    logic s1219 ,c1219; 
    fa fa1219 (pp_25_59, pp_26_57, pp_27_55, s1219, c1219);
    logic s1220 ,c1220; 
    fa fa1220 (const1, pp_23_64, pp_24_62, s1220, c1220);
    logic s1221 ,c1221;
    ha ha1221 (pp_25_60, pp_26_58, s1221, c1221);
    logic s1222 ,c1222; 
    fa fa1222 (pp_23_65, pp_24_63, pp_25_61, s1222, c1222);
    logic s1223 ,c1223;
    ha ha1223 (const1, pp_24_64, s1223, c1223);
    logic s1224 ,c1224;
    ha ha1224 (pp_0_10, pp_1_8, s1224, c1224);
    logic s1225 ,c1225;
    ha ha1225 (pp_0_11, pp_1_9, s1225, c1225);
    logic s1226 ,c1226; 
    fa fa1226 (pp_0_12, pp_1_10, pp_2_8, s1226, c1226);
    logic s1227 ,c1227;
    ha ha1227 (pp_3_6, pp_4_4, s1227, c1227);
    logic s1228 ,c1228; 
    fa fa1228 (pp_0_13, pp_1_11, pp_2_9, s1228, c1228);
    logic s1229 ,c1229;
    ha ha1229 (pp_3_7, pp_4_5, s1229, c1229);
    logic s1230 ,c1230; 
    fa fa1230 (pp_0_14, pp_1_12, pp_2_10, s1230, c1230);
    logic s1231 ,c1231; 
    fa fa1231 (pp_3_8, pp_4_6, pp_5_4, s1231, c1231);
    logic s1232 ,c1232;
    ha ha1232 (pp_6_2, pp_7_0, s1232, c1232);
    logic s1233 ,c1233; 
    fa fa1233 (pp_0_15, pp_1_13, pp_2_11, s1233, c1233);
    logic s1234 ,c1234; 
    fa fa1234 (pp_3_9, pp_4_7, pp_5_5, s1234, c1234);
    logic s1235 ,c1235;
    ha ha1235 (pp_6_3, pp_7_1, s1235, c1235);
    logic s1236 ,c1236; 
    fa fa1236 (pp_2_12, pp_3_10, pp_4_8, s1236, c1236);
    logic s1237 ,c1237; 
    fa fa1237 (pp_5_6, pp_6_4, pp_7_2, s1237, c1237);
    logic s1238 ,c1238; 
    fa fa1238 (pp_8_0, tcomp8, s860, s1238, c1238);
    logic s1239 ,c1239; 
    fa fa1239 (pp_2_13, pp_3_11, pp_4_9, s1239, c1239);
    logic s1240 ,c1240; 
    fa fa1240 (pp_5_7, pp_6_5, pp_7_3, s1240, c1240);
    logic s1241 ,c1241; 
    fa fa1241 (pp_8_1, c860, s861, s1241, c1241);
    logic s1242 ,c1242; 
    fa fa1242 (pp_5_8, pp_6_6, pp_7_4, s1242, c1242);
    logic s1243 ,c1243; 
    fa fa1243 (pp_8_2, pp_9_0, tcomp9, s1243, c1243);
    logic s1244 ,c1244; 
    fa fa1244 (c861, s862, s863, s1244, c1244);
    logic s1245 ,c1245; 
    fa fa1245 (pp_5_9, pp_6_7, pp_7_5, s1245, c1245);
    logic s1246 ,c1246; 
    fa fa1246 (pp_8_3, pp_9_1, c862, s1246, c1246);
    logic s1247 ,c1247; 
    fa fa1247 (c863, s864, s865, s1247, c1247);
    logic s1248 ,c1248; 
    fa fa1248 (pp_8_4, pp_9_2, pp_10_0, s1248, c1248);
    logic s1249 ,c1249; 
    fa fa1249 (tcomp10, c864, c865, s1249, c1249);
    logic s1250 ,c1250; 
    fa fa1250 (s866, s867, s868, s1250, c1250);
    logic s1251 ,c1251; 
    fa fa1251 (pp_8_5, pp_9_3, pp_10_1, s1251, c1251);
    logic s1252 ,c1252; 
    fa fa1252 (c866, c867, c868, s1252, c1252);
    logic s1253 ,c1253; 
    fa fa1253 (s869, s870, s871, s1253, c1253);
    logic s1254 ,c1254; 
    fa fa1254 (pp_11_0, tcomp11, c869, s1254, c1254);
    logic s1255 ,c1255; 
    fa fa1255 (c870, c871, s872, s1255, c1255);
    logic s1256 ,c1256; 
    fa fa1256 (s873, s874, s875, s1256, c1256);
    logic s1257 ,c1257; 
    fa fa1257 (pp_11_1, c872, c873, s1257, c1257);
    logic s1258 ,c1258; 
    fa fa1258 (c874, c875, s876, s1258, c1258);
    logic s1259 ,c1259; 
    fa fa1259 (s877, s878, s879, s1259, c1259);
    logic s1260 ,c1260; 
    fa fa1260 (s434, c876, c877, s1260, c1260);
    logic s1261 ,c1261; 
    fa fa1261 (c878, c879, s880, s1261, c1261);
    logic s1262 ,c1262; 
    fa fa1262 (s881, s882, s883, s1262, c1262);
    logic s1263 ,c1263; 
    fa fa1263 (s435, c880, c881, s1263, c1263);
    logic s1264 ,c1264; 
    fa fa1264 (c882, c883, s884, s1264, c1264);
    logic s1265 ,c1265; 
    fa fa1265 (s885, s886, s887, s1265, c1265);
    logic s1266 ,c1266; 
    fa fa1266 (s437, c884, c885, s1266, c1266);
    logic s1267 ,c1267; 
    fa fa1267 (c886, c887, s888, s1267, c1267);
    logic s1268 ,c1268; 
    fa fa1268 (s889, s890, s891, s1268, c1268);
    logic s1269 ,c1269; 
    fa fa1269 (s439, c888, c889, s1269, c1269);
    logic s1270 ,c1270; 
    fa fa1270 (c890, c891, s892, s1270, c1270);
    logic s1271 ,c1271; 
    fa fa1271 (s893, s894, s895, s1271, c1271);
    logic s1272 ,c1272; 
    fa fa1272 (s442, c892, c893, s1272, c1272);
    logic s1273 ,c1273; 
    fa fa1273 (c894, c895, s896, s1273, c1273);
    logic s1274 ,c1274; 
    fa fa1274 (s897, s898, s899, s1274, c1274);
    logic s1275 ,c1275; 
    fa fa1275 (s445, c896, c897, s1275, c1275);
    logic s1276 ,c1276; 
    fa fa1276 (c898, c899, s900, s1276, c1276);
    logic s1277 ,c1277; 
    fa fa1277 (s901, s902, s903, s1277, c1277);
    logic s1278 ,c1278; 
    fa fa1278 (s449, c900, c901, s1278, c1278);
    logic s1279 ,c1279; 
    fa fa1279 (c902, c903, s904, s1279, c1279);
    logic s1280 ,c1280; 
    fa fa1280 (s905, s906, s907, s1280, c1280);
    logic s1281 ,c1281; 
    fa fa1281 (s453, c904, c905, s1281, c1281);
    logic s1282 ,c1282; 
    fa fa1282 (c906, c907, s908, s1282, c1282);
    logic s1283 ,c1283; 
    fa fa1283 (s909, s910, s911, s1283, c1283);
    logic s1284 ,c1284; 
    fa fa1284 (s458, c908, c909, s1284, c1284);
    logic s1285 ,c1285; 
    fa fa1285 (c910, c911, s912, s1285, c1285);
    logic s1286 ,c1286; 
    fa fa1286 (s913, s914, s915, s1286, c1286);
    logic s1287 ,c1287; 
    fa fa1287 (s463, c912, c913, s1287, c1287);
    logic s1288 ,c1288; 
    fa fa1288 (c914, c915, s916, s1288, c1288);
    logic s1289 ,c1289; 
    fa fa1289 (s917, s918, s919, s1289, c1289);
    logic s1290 ,c1290; 
    fa fa1290 (s469, c916, c917, s1290, c1290);
    logic s1291 ,c1291; 
    fa fa1291 (c918, c919, s920, s1291, c1291);
    logic s1292 ,c1292; 
    fa fa1292 (s921, s922, s923, s1292, c1292);
    logic s1293 ,c1293; 
    fa fa1293 (s475, c920, c921, s1293, c1293);
    logic s1294 ,c1294; 
    fa fa1294 (c922, c923, s924, s1294, c1294);
    logic s1295 ,c1295; 
    fa fa1295 (s925, s926, s927, s1295, c1295);
    logic s1296 ,c1296; 
    fa fa1296 (s481, c924, c925, s1296, c1296);
    logic s1297 ,c1297; 
    fa fa1297 (c926, c927, s928, s1297, c1297);
    logic s1298 ,c1298; 
    fa fa1298 (s929, s930, s931, s1298, c1298);
    logic s1299 ,c1299; 
    fa fa1299 (s487, c928, c929, s1299, c1299);
    logic s1300 ,c1300; 
    fa fa1300 (c930, c931, s932, s1300, c1300);
    logic s1301 ,c1301; 
    fa fa1301 (s933, s934, s935, s1301, c1301);
    logic s1302 ,c1302; 
    fa fa1302 (s493, c932, c933, s1302, c1302);
    logic s1303 ,c1303; 
    fa fa1303 (c934, c935, s936, s1303, c1303);
    logic s1304 ,c1304; 
    fa fa1304 (s937, s938, s939, s1304, c1304);
    logic s1305 ,c1305; 
    fa fa1305 (s499, c936, c937, s1305, c1305);
    logic s1306 ,c1306; 
    fa fa1306 (c938, c939, s940, s1306, c1306);
    logic s1307 ,c1307; 
    fa fa1307 (s941, s942, s943, s1307, c1307);
    logic s1308 ,c1308; 
    fa fa1308 (s505, c940, c941, s1308, c1308);
    logic s1309 ,c1309; 
    fa fa1309 (c942, c943, s944, s1309, c1309);
    logic s1310 ,c1310; 
    fa fa1310 (s945, s946, s947, s1310, c1310);
    logic s1311 ,c1311; 
    fa fa1311 (s511, c944, c945, s1311, c1311);
    logic s1312 ,c1312; 
    fa fa1312 (c946, c947, s948, s1312, c1312);
    logic s1313 ,c1313; 
    fa fa1313 (s949, s950, s951, s1313, c1313);
    logic s1314 ,c1314; 
    fa fa1314 (s517, c948, c949, s1314, c1314);
    logic s1315 ,c1315; 
    fa fa1315 (c950, c951, s952, s1315, c1315);
    logic s1316 ,c1316; 
    fa fa1316 (s953, s954, s955, s1316, c1316);
    logic s1317 ,c1317; 
    fa fa1317 (s523, c952, c953, s1317, c1317);
    logic s1318 ,c1318; 
    fa fa1318 (c954, c955, s956, s1318, c1318);
    logic s1319 ,c1319; 
    fa fa1319 (s957, s958, s959, s1319, c1319);
    logic s1320 ,c1320; 
    fa fa1320 (s529, c956, c957, s1320, c1320);
    logic s1321 ,c1321; 
    fa fa1321 (c958, c959, s960, s1321, c1321);
    logic s1322 ,c1322; 
    fa fa1322 (s961, s962, s963, s1322, c1322);
    logic s1323 ,c1323; 
    fa fa1323 (s535, c960, c961, s1323, c1323);
    logic s1324 ,c1324; 
    fa fa1324 (c962, c963, s964, s1324, c1324);
    logic s1325 ,c1325; 
    fa fa1325 (s965, s966, s967, s1325, c1325);
    logic s1326 ,c1326; 
    fa fa1326 (s541, c964, c965, s1326, c1326);
    logic s1327 ,c1327; 
    fa fa1327 (c966, c967, s968, s1327, c1327);
    logic s1328 ,c1328; 
    fa fa1328 (s969, s970, s971, s1328, c1328);
    logic s1329 ,c1329; 
    fa fa1329 (s547, c968, c969, s1329, c1329);
    logic s1330 ,c1330; 
    fa fa1330 (c970, c971, s972, s1330, c1330);
    logic s1331 ,c1331; 
    fa fa1331 (s973, s974, s975, s1331, c1331);
    logic s1332 ,c1332; 
    fa fa1332 (s553, c972, c973, s1332, c1332);
    logic s1333 ,c1333; 
    fa fa1333 (c974, c975, s976, s1333, c1333);
    logic s1334 ,c1334; 
    fa fa1334 (s977, s978, s979, s1334, c1334);
    logic s1335 ,c1335; 
    fa fa1335 (s559, c976, c977, s1335, c1335);
    logic s1336 ,c1336; 
    fa fa1336 (c978, c979, s980, s1336, c1336);
    logic s1337 ,c1337; 
    fa fa1337 (s981, s982, s983, s1337, c1337);
    logic s1338 ,c1338; 
    fa fa1338 (s565, c980, c981, s1338, c1338);
    logic s1339 ,c1339; 
    fa fa1339 (c982, c983, s984, s1339, c1339);
    logic s1340 ,c1340; 
    fa fa1340 (s985, s986, s987, s1340, c1340);
    logic s1341 ,c1341; 
    fa fa1341 (s571, c984, c985, s1341, c1341);
    logic s1342 ,c1342; 
    fa fa1342 (c986, c987, s988, s1342, c1342);
    logic s1343 ,c1343; 
    fa fa1343 (s989, s990, s991, s1343, c1343);
    logic s1344 ,c1344; 
    fa fa1344 (s577, c988, c989, s1344, c1344);
    logic s1345 ,c1345; 
    fa fa1345 (c990, c991, s992, s1345, c1345);
    logic s1346 ,c1346; 
    fa fa1346 (s993, s994, s995, s1346, c1346);
    logic s1347 ,c1347; 
    fa fa1347 (s583, c992, c993, s1347, c1347);
    logic s1348 ,c1348; 
    fa fa1348 (c994, c995, s996, s1348, c1348);
    logic s1349 ,c1349; 
    fa fa1349 (s997, s998, s999, s1349, c1349);
    logic s1350 ,c1350; 
    fa fa1350 (s589, c996, c997, s1350, c1350);
    logic s1351 ,c1351; 
    fa fa1351 (c998, c999, s1000, s1351, c1351);
    logic s1352 ,c1352; 
    fa fa1352 (s1001, s1002, s1003, s1352, c1352);
    logic s1353 ,c1353; 
    fa fa1353 (s595, c1000, c1001, s1353, c1353);
    logic s1354 ,c1354; 
    fa fa1354 (c1002, c1003, s1004, s1354, c1354);
    logic s1355 ,c1355; 
    fa fa1355 (s1005, s1006, s1007, s1355, c1355);
    logic s1356 ,c1356; 
    fa fa1356 (s601, c1004, c1005, s1356, c1356);
    logic s1357 ,c1357; 
    fa fa1357 (c1006, c1007, s1008, s1357, c1357);
    logic s1358 ,c1358; 
    fa fa1358 (s1009, s1010, s1011, s1358, c1358);
    logic s1359 ,c1359; 
    fa fa1359 (s607, c1008, c1009, s1359, c1359);
    logic s1360 ,c1360; 
    fa fa1360 (c1010, c1011, s1012, s1360, c1360);
    logic s1361 ,c1361; 
    fa fa1361 (s1013, s1014, s1015, s1361, c1361);
    logic s1362 ,c1362; 
    fa fa1362 (s613, c1012, c1013, s1362, c1362);
    logic s1363 ,c1363; 
    fa fa1363 (c1014, c1015, s1016, s1363, c1363);
    logic s1364 ,c1364; 
    fa fa1364 (s1017, s1018, s1019, s1364, c1364);
    logic s1365 ,c1365; 
    fa fa1365 (s619, c1016, c1017, s1365, c1365);
    logic s1366 ,c1366; 
    fa fa1366 (c1018, c1019, s1020, s1366, c1366);
    logic s1367 ,c1367; 
    fa fa1367 (s1021, s1022, s1023, s1367, c1367);
    logic s1368 ,c1368; 
    fa fa1368 (s625, c1020, c1021, s1368, c1368);
    logic s1369 ,c1369; 
    fa fa1369 (c1022, c1023, s1024, s1369, c1369);
    logic s1370 ,c1370; 
    fa fa1370 (s1025, s1026, s1027, s1370, c1370);
    logic s1371 ,c1371; 
    fa fa1371 (s631, c1024, c1025, s1371, c1371);
    logic s1372 ,c1372; 
    fa fa1372 (c1026, c1027, s1028, s1372, c1372);
    logic s1373 ,c1373; 
    fa fa1373 (s1029, s1030, s1031, s1373, c1373);
    logic s1374 ,c1374; 
    fa fa1374 (s637, c1028, c1029, s1374, c1374);
    logic s1375 ,c1375; 
    fa fa1375 (c1030, c1031, s1032, s1375, c1375);
    logic s1376 ,c1376; 
    fa fa1376 (s1033, s1034, s1035, s1376, c1376);
    logic s1377 ,c1377; 
    fa fa1377 (s643, c1032, c1033, s1377, c1377);
    logic s1378 ,c1378; 
    fa fa1378 (c1034, c1035, s1036, s1378, c1378);
    logic s1379 ,c1379; 
    fa fa1379 (s1037, s1038, s1039, s1379, c1379);
    logic s1380 ,c1380; 
    fa fa1380 (s649, c1036, c1037, s1380, c1380);
    logic s1381 ,c1381; 
    fa fa1381 (c1038, c1039, s1040, s1381, c1381);
    logic s1382 ,c1382; 
    fa fa1382 (s1041, s1042, s1043, s1382, c1382);
    logic s1383 ,c1383; 
    fa fa1383 (s655, c1040, c1041, s1383, c1383);
    logic s1384 ,c1384; 
    fa fa1384 (c1042, c1043, s1044, s1384, c1384);
    logic s1385 ,c1385; 
    fa fa1385 (s1045, s1046, s1047, s1385, c1385);
    logic s1386 ,c1386; 
    fa fa1386 (s661, c1044, c1045, s1386, c1386);
    logic s1387 ,c1387; 
    fa fa1387 (c1046, c1047, s1048, s1387, c1387);
    logic s1388 ,c1388; 
    fa fa1388 (s1049, s1050, s1051, s1388, c1388);
    logic s1389 ,c1389; 
    fa fa1389 (s667, c1048, c1049, s1389, c1389);
    logic s1390 ,c1390; 
    fa fa1390 (c1050, c1051, s1052, s1390, c1390);
    logic s1391 ,c1391; 
    fa fa1391 (s1053, s1054, s1055, s1391, c1391);
    logic s1392 ,c1392; 
    fa fa1392 (s673, c1052, c1053, s1392, c1392);
    logic s1393 ,c1393; 
    fa fa1393 (c1054, c1055, s1056, s1393, c1393);
    logic s1394 ,c1394; 
    fa fa1394 (s1057, s1058, s1059, s1394, c1394);
    logic s1395 ,c1395; 
    fa fa1395 (s679, c1056, c1057, s1395, c1395);
    logic s1396 ,c1396; 
    fa fa1396 (c1058, c1059, s1060, s1396, c1396);
    logic s1397 ,c1397; 
    fa fa1397 (s1061, s1062, s1063, s1397, c1397);
    logic s1398 ,c1398; 
    fa fa1398 (s685, c1060, c1061, s1398, c1398);
    logic s1399 ,c1399; 
    fa fa1399 (c1062, c1063, s1064, s1399, c1399);
    logic s1400 ,c1400; 
    fa fa1400 (s1065, s1066, s1067, s1400, c1400);
    logic s1401 ,c1401; 
    fa fa1401 (s691, c1064, c1065, s1401, c1401);
    logic s1402 ,c1402; 
    fa fa1402 (c1066, c1067, s1068, s1402, c1402);
    logic s1403 ,c1403; 
    fa fa1403 (s1069, s1070, s1071, s1403, c1403);
    logic s1404 ,c1404; 
    fa fa1404 (s697, c1068, c1069, s1404, c1404);
    logic s1405 ,c1405; 
    fa fa1405 (c1070, c1071, s1072, s1405, c1405);
    logic s1406 ,c1406; 
    fa fa1406 (s1073, s1074, s1075, s1406, c1406);
    logic s1407 ,c1407; 
    fa fa1407 (s703, c1072, c1073, s1407, c1407);
    logic s1408 ,c1408; 
    fa fa1408 (c1074, c1075, s1076, s1408, c1408);
    logic s1409 ,c1409; 
    fa fa1409 (s1077, s1078, s1079, s1409, c1409);
    logic s1410 ,c1410; 
    fa fa1410 (s709, c1076, c1077, s1410, c1410);
    logic s1411 ,c1411; 
    fa fa1411 (c1078, c1079, s1080, s1411, c1411);
    logic s1412 ,c1412; 
    fa fa1412 (s1081, s1082, s1083, s1412, c1412);
    logic s1413 ,c1413; 
    fa fa1413 (s715, c1080, c1081, s1413, c1413);
    logic s1414 ,c1414; 
    fa fa1414 (c1082, c1083, s1084, s1414, c1414);
    logic s1415 ,c1415; 
    fa fa1415 (s1085, s1086, s1087, s1415, c1415);
    logic s1416 ,c1416; 
    fa fa1416 (s721, c1084, c1085, s1416, c1416);
    logic s1417 ,c1417; 
    fa fa1417 (c1086, c1087, s1088, s1417, c1417);
    logic s1418 ,c1418; 
    fa fa1418 (s1089, s1090, s1091, s1418, c1418);
    logic s1419 ,c1419; 
    fa fa1419 (s727, c1088, c1089, s1419, c1419);
    logic s1420 ,c1420; 
    fa fa1420 (c1090, c1091, s1092, s1420, c1420);
    logic s1421 ,c1421; 
    fa fa1421 (s1093, s1094, s1095, s1421, c1421);
    logic s1422 ,c1422; 
    fa fa1422 (s733, c1092, c1093, s1422, c1422);
    logic s1423 ,c1423; 
    fa fa1423 (c1094, c1095, s1096, s1423, c1423);
    logic s1424 ,c1424; 
    fa fa1424 (s1097, s1098, s1099, s1424, c1424);
    logic s1425 ,c1425; 
    fa fa1425 (s739, c1096, c1097, s1425, c1425);
    logic s1426 ,c1426; 
    fa fa1426 (c1098, c1099, s1100, s1426, c1426);
    logic s1427 ,c1427; 
    fa fa1427 (s1101, s1102, s1103, s1427, c1427);
    logic s1428 ,c1428; 
    fa fa1428 (s745, c1100, c1101, s1428, c1428);
    logic s1429 ,c1429; 
    fa fa1429 (c1102, c1103, s1104, s1429, c1429);
    logic s1430 ,c1430; 
    fa fa1430 (s1105, s1106, s1107, s1430, c1430);
    logic s1431 ,c1431; 
    fa fa1431 (s751, c1104, c1105, s1431, c1431);
    logic s1432 ,c1432; 
    fa fa1432 (c1106, c1107, s1108, s1432, c1432);
    logic s1433 ,c1433; 
    fa fa1433 (s1109, s1110, s1111, s1433, c1433);
    logic s1434 ,c1434; 
    fa fa1434 (s757, c1108, c1109, s1434, c1434);
    logic s1435 ,c1435; 
    fa fa1435 (c1110, c1111, s1112, s1435, c1435);
    logic s1436 ,c1436; 
    fa fa1436 (s1113, s1114, s1115, s1436, c1436);
    logic s1437 ,c1437; 
    fa fa1437 (s763, c1112, c1113, s1437, c1437);
    logic s1438 ,c1438; 
    fa fa1438 (c1114, c1115, s1116, s1438, c1438);
    logic s1439 ,c1439; 
    fa fa1439 (s1117, s1118, s1119, s1439, c1439);
    logic s1440 ,c1440; 
    fa fa1440 (s769, c1116, c1117, s1440, c1440);
    logic s1441 ,c1441; 
    fa fa1441 (c1118, c1119, s1120, s1441, c1441);
    logic s1442 ,c1442; 
    fa fa1442 (s1121, s1122, s1123, s1442, c1442);
    logic s1443 ,c1443; 
    fa fa1443 (s775, c1120, c1121, s1443, c1443);
    logic s1444 ,c1444; 
    fa fa1444 (c1122, c1123, s1124, s1444, c1444);
    logic s1445 ,c1445; 
    fa fa1445 (s1125, s1126, s1127, s1445, c1445);
    logic s1446 ,c1446; 
    fa fa1446 (s781, c1124, c1125, s1446, c1446);
    logic s1447 ,c1447; 
    fa fa1447 (c1126, c1127, s1128, s1447, c1447);
    logic s1448 ,c1448; 
    fa fa1448 (s1129, s1130, s1131, s1448, c1448);
    logic s1449 ,c1449; 
    fa fa1449 (s787, c1128, c1129, s1449, c1449);
    logic s1450 ,c1450; 
    fa fa1450 (c1130, c1131, s1132, s1450, c1450);
    logic s1451 ,c1451; 
    fa fa1451 (s1133, s1134, s1135, s1451, c1451);
    logic s1452 ,c1452; 
    fa fa1452 (s793, c1132, c1133, s1452, c1452);
    logic s1453 ,c1453; 
    fa fa1453 (c1134, c1135, s1136, s1453, c1453);
    logic s1454 ,c1454; 
    fa fa1454 (s1137, s1138, s1139, s1454, c1454);
    logic s1455 ,c1455; 
    fa fa1455 (s799, c1136, c1137, s1455, c1455);
    logic s1456 ,c1456; 
    fa fa1456 (c1138, c1139, s1140, s1456, c1456);
    logic s1457 ,c1457; 
    fa fa1457 (s1141, s1142, s1143, s1457, c1457);
    logic s1458 ,c1458; 
    fa fa1458 (s805, c1140, c1141, s1458, c1458);
    logic s1459 ,c1459; 
    fa fa1459 (c1142, c1143, s1144, s1459, c1459);
    logic s1460 ,c1460; 
    fa fa1460 (s1145, s1146, s1147, s1460, c1460);
    logic s1461 ,c1461; 
    fa fa1461 (s811, c1144, c1145, s1461, c1461);
    logic s1462 ,c1462; 
    fa fa1462 (c1146, c1147, s1148, s1462, c1462);
    logic s1463 ,c1463; 
    fa fa1463 (s1149, s1150, s1151, s1463, c1463);
    logic s1464 ,c1464; 
    fa fa1464 (s817, c1148, c1149, s1464, c1464);
    logic s1465 ,c1465; 
    fa fa1465 (c1150, c1151, s1152, s1465, c1465);
    logic s1466 ,c1466; 
    fa fa1466 (s1153, s1154, s1155, s1466, c1466);
    logic s1467 ,c1467; 
    fa fa1467 (s823, c1152, c1153, s1467, c1467);
    logic s1468 ,c1468; 
    fa fa1468 (c1154, c1155, s1156, s1468, c1468);
    logic s1469 ,c1469; 
    fa fa1469 (s1157, s1158, s1159, s1469, c1469);
    logic s1470 ,c1470; 
    fa fa1470 (s829, c1156, c1157, s1470, c1470);
    logic s1471 ,c1471; 
    fa fa1471 (c1158, c1159, s1160, s1471, c1471);
    logic s1472 ,c1472; 
    fa fa1472 (s1161, s1162, s1163, s1472, c1472);
    logic s1473 ,c1473; 
    fa fa1473 (s834, c1160, c1161, s1473, c1473);
    logic s1474 ,c1474; 
    fa fa1474 (c1162, c1163, s1164, s1474, c1474);
    logic s1475 ,c1475; 
    fa fa1475 (s1165, s1166, s1167, s1475, c1475);
    logic s1476 ,c1476; 
    fa fa1476 (s839, c1164, c1165, s1476, c1476);
    logic s1477 ,c1477; 
    fa fa1477 (c1166, c1167, s1168, s1477, c1477);
    logic s1478 ,c1478; 
    fa fa1478 (s1169, s1170, s1171, s1478, c1478);
    logic s1479 ,c1479; 
    fa fa1479 (s843, c1168, c1169, s1479, c1479);
    logic s1480 ,c1480; 
    fa fa1480 (c1170, c1171, s1172, s1480, c1480);
    logic s1481 ,c1481; 
    fa fa1481 (s1173, s1174, s1175, s1481, c1481);
    logic s1482 ,c1482; 
    fa fa1482 (s847, c1172, c1173, s1482, c1482);
    logic s1483 ,c1483; 
    fa fa1483 (c1174, c1175, s1176, s1483, c1483);
    logic s1484 ,c1484; 
    fa fa1484 (s1177, s1178, s1179, s1484, c1484);
    logic s1485 ,c1485; 
    fa fa1485 (s850, c1176, c1177, s1485, c1485);
    logic s1486 ,c1486; 
    fa fa1486 (c1178, c1179, s1180, s1486, c1486);
    logic s1487 ,c1487; 
    fa fa1487 (s1181, s1182, s1183, s1487, c1487);
    logic s1488 ,c1488; 
    fa fa1488 (s853, c1180, c1181, s1488, c1488);
    logic s1489 ,c1489; 
    fa fa1489 (c1182, c1183, s1184, s1489, c1489);
    logic s1490 ,c1490; 
    fa fa1490 (s1185, s1186, s1187, s1490, c1490);
    logic s1491 ,c1491; 
    fa fa1491 (s855, c1184, c1185, s1491, c1491);
    logic s1492 ,c1492; 
    fa fa1492 (c1186, c1187, s1188, s1492, c1492);
    logic s1493 ,c1493; 
    fa fa1493 (s1189, s1190, s1191, s1493, c1493);
    logic s1494 ,c1494; 
    fa fa1494 (s857, c1188, c1189, s1494, c1494);
    logic s1495 ,c1495; 
    fa fa1495 (c1190, c1191, s1192, s1495, c1495);
    logic s1496 ,c1496; 
    fa fa1496 (s1193, s1194, s1195, s1496, c1496);
    logic s1497 ,c1497; 
    fa fa1497 (s858, c1192, c1193, s1497, c1497);
    logic s1498 ,c1498; 
    fa fa1498 (c1194, c1195, s1196, s1498, c1498);
    logic s1499 ,c1499; 
    fa fa1499 (s1197, s1198, s1199, s1499, c1499);
    logic s1500 ,c1500; 
    fa fa1500 (s859, c1196, c1197, s1500, c1500);
    logic s1501 ,c1501; 
    fa fa1501 (c1198, c1199, s1200, s1501, c1501);
    logic s1502 ,c1502; 
    fa fa1502 (s1201, s1202, s1203, s1502, c1502);
    logic s1503 ,c1503; 
    fa fa1503 (c859, c1200, c1201, s1503, c1503);
    logic s1504 ,c1504; 
    fa fa1504 (c1202, c1203, s1204, s1504, c1504);
    logic s1505 ,c1505; 
    fa fa1505 (s1205, s1206, s1207, s1505, c1505);
    logic s1506 ,c1506; 
    fa fa1506 (pp_31_44, c1204, c1205, s1506, c1506);
    logic s1507 ,c1507; 
    fa fa1507 (c1206, c1207, s1208, s1507, c1507);
    logic s1508 ,c1508; 
    fa fa1508 (s1209, s1210, s1211, s1508, c1508);
    logic s1509 ,c1509; 
    fa fa1509 (pp_30_47, pp_31_45, c1208, s1509, c1509);
    logic s1510 ,c1510; 
    fa fa1510 (c1209, c1210, c1211, s1510, c1510);
    logic s1511 ,c1511; 
    fa fa1511 (s1212, s1213, s1214, s1511, c1511);
    logic s1512 ,c1512; 
    fa fa1512 (pp_29_50, pp_30_48, pp_31_46, s1512, c1512);
    logic s1513 ,c1513; 
    fa fa1513 (c1212, c1213, c1214, s1513, c1513);
    logic s1514 ,c1514; 
    fa fa1514 (s1215, s1216, s1217, s1514, c1514);
    logic s1515 ,c1515; 
    fa fa1515 (pp_28_53, pp_29_51, pp_30_49, s1515, c1515);
    logic s1516 ,c1516; 
    fa fa1516 (pp_31_47, c1215, c1216, s1516, c1516);
    logic s1517 ,c1517; 
    fa fa1517 (c1217, s1218, s1219, s1517, c1517);
    logic s1518 ,c1518; 
    fa fa1518 (pp_27_56, pp_28_54, pp_29_52, s1518, c1518);
    logic s1519 ,c1519; 
    fa fa1519 (pp_30_50, pp_31_48, c1218, s1519, c1519);
    logic s1520 ,c1520; 
    fa fa1520 (c1219, s1220, s1221, s1520, c1520);
    logic s1521 ,c1521; 
    fa fa1521 (pp_26_59, pp_27_57, pp_28_55, s1521, c1521);
    logic s1522 ,c1522; 
    fa fa1522 (pp_29_53, pp_30_51, pp_31_49, s1522, c1522);
    logic s1523 ,c1523; 
    fa fa1523 (c1220, c1221, s1222, s1523, c1523);
    logic s1524 ,c1524; 
    fa fa1524 (pp_25_62, pp_26_60, pp_27_58, s1524, c1524);
    logic s1525 ,c1525; 
    fa fa1525 (pp_28_56, pp_29_54, pp_30_52, s1525, c1525);
    logic s1526 ,c1526; 
    fa fa1526 (pp_31_50, c1222, s1223, s1526, c1526);
    logic s1527 ,c1527; 
    fa fa1527 (pp_24_65, pp_25_63, pp_26_61, s1527, c1527);
    logic s1528 ,c1528; 
    fa fa1528 (pp_27_59, pp_28_57, pp_29_55, s1528, c1528);
    logic s1529 ,c1529; 
    fa fa1529 (pp_30_53, pp_31_51, c1223, s1529, c1529);
    logic s1530 ,c1530; 
    fa fa1530 (const1, pp_25_64, pp_26_62, s1530, c1530);
    logic s1531 ,c1531; 
    fa fa1531 (pp_27_60, pp_28_58, pp_29_56, s1531, c1531);
    logic s1532 ,c1532;
    ha ha1532 (pp_30_54, pp_31_52, s1532, c1532);
    logic s1533 ,c1533; 
    fa fa1533 (pp_25_65, pp_26_63, pp_27_61, s1533, c1533);
    logic s1534 ,c1534; 
    fa fa1534 (pp_28_59, pp_29_57, pp_30_55, s1534, c1534);
    logic s1535 ,c1535; 
    fa fa1535 (const1, pp_26_64, pp_27_62, s1535, c1535);
    logic s1536 ,c1536;
    ha ha1536 (pp_28_60, pp_29_58, s1536, c1536);
    logic s1537 ,c1537; 
    fa fa1537 (pp_26_65, pp_27_63, pp_28_61, s1537, c1537);
    logic s1538 ,c1538;
    ha ha1538 (const1, pp_27_64, s1538, c1538);
    logic s1539 ,c1539;
    ha ha1539 (pp_0_6, pp_1_4, s1539, c1539);
    logic s1540 ,c1540;
    ha ha1540 (pp_0_7, pp_1_5, s1540, c1540);
    logic s1541 ,c1541; 
    fa fa1541 (pp_0_8, pp_1_6, pp_2_4, s1541, c1541);
    logic s1542 ,c1542;
    ha ha1542 (pp_3_2, pp_4_0, s1542, c1542);
    logic s1543 ,c1543; 
    fa fa1543 (pp_0_9, pp_1_7, pp_2_5, s1543, c1543);
    logic s1544 ,c1544;
    ha ha1544 (pp_3_3, pp_4_1, s1544, c1544);
    logic s1545 ,c1545; 
    fa fa1545 (pp_2_6, pp_3_4, pp_4_2, s1545, c1545);
    logic s1546 ,c1546; 
    fa fa1546 (pp_5_0, tcomp5, s1224, s1546, c1546);
    logic s1547 ,c1547; 
    fa fa1547 (pp_2_7, pp_3_5, pp_4_3, s1547, c1547);
    logic s1548 ,c1548; 
    fa fa1548 (pp_5_1, c1224, s1225, s1548, c1548);
    logic s1549 ,c1549; 
    fa fa1549 (pp_5_2, pp_6_0, tcomp6, s1549, c1549);
    logic s1550 ,c1550; 
    fa fa1550 (c1225, s1226, s1227, s1550, c1550);
    logic s1551 ,c1551; 
    fa fa1551 (pp_5_3, pp_6_1, c1226, s1551, c1551);
    logic s1552 ,c1552; 
    fa fa1552 (c1227, s1228, s1229, s1552, c1552);
    logic s1553 ,c1553; 
    fa fa1553 (tcomp7, c1228, c1229, s1553, c1553);
    logic s1554 ,c1554; 
    fa fa1554 (s1230, s1231, s1232, s1554, c1554);
    logic s1555 ,c1555; 
    fa fa1555 (c1230, c1231, c1232, s1555, c1555);
    logic s1556 ,c1556; 
    fa fa1556 (s1233, s1234, s1235, s1556, c1556);
    logic s1557 ,c1557; 
    fa fa1557 (c1233, c1234, c1235, s1557, c1557);
    logic s1558 ,c1558; 
    fa fa1558 (s1236, s1237, s1238, s1558, c1558);
    logic s1559 ,c1559; 
    fa fa1559 (c1236, c1237, c1238, s1559, c1559);
    logic s1560 ,c1560; 
    fa fa1560 (s1239, s1240, s1241, s1560, c1560);
    logic s1561 ,c1561; 
    fa fa1561 (c1239, c1240, c1241, s1561, c1561);
    logic s1562 ,c1562; 
    fa fa1562 (s1242, s1243, s1244, s1562, c1562);
    logic s1563 ,c1563; 
    fa fa1563 (c1242, c1243, c1244, s1563, c1563);
    logic s1564 ,c1564; 
    fa fa1564 (s1245, s1246, s1247, s1564, c1564);
    logic s1565 ,c1565; 
    fa fa1565 (c1245, c1246, c1247, s1565, c1565);
    logic s1566 ,c1566; 
    fa fa1566 (s1248, s1249, s1250, s1566, c1566);
    logic s1567 ,c1567; 
    fa fa1567 (c1248, c1249, c1250, s1567, c1567);
    logic s1568 ,c1568; 
    fa fa1568 (s1251, s1252, s1253, s1568, c1568);
    logic s1569 ,c1569; 
    fa fa1569 (c1251, c1252, c1253, s1569, c1569);
    logic s1570 ,c1570; 
    fa fa1570 (s1254, s1255, s1256, s1570, c1570);
    logic s1571 ,c1571; 
    fa fa1571 (c1254, c1255, c1256, s1571, c1571);
    logic s1572 ,c1572; 
    fa fa1572 (s1257, s1258, s1259, s1572, c1572);
    logic s1573 ,c1573; 
    fa fa1573 (c1257, c1258, c1259, s1573, c1573);
    logic s1574 ,c1574; 
    fa fa1574 (s1260, s1261, s1262, s1574, c1574);
    logic s1575 ,c1575; 
    fa fa1575 (c1260, c1261, c1262, s1575, c1575);
    logic s1576 ,c1576; 
    fa fa1576 (s1263, s1264, s1265, s1576, c1576);
    logic s1577 ,c1577; 
    fa fa1577 (c1263, c1264, c1265, s1577, c1577);
    logic s1578 ,c1578; 
    fa fa1578 (s1266, s1267, s1268, s1578, c1578);
    logic s1579 ,c1579; 
    fa fa1579 (c1266, c1267, c1268, s1579, c1579);
    logic s1580 ,c1580; 
    fa fa1580 (s1269, s1270, s1271, s1580, c1580);
    logic s1581 ,c1581; 
    fa fa1581 (c1269, c1270, c1271, s1581, c1581);
    logic s1582 ,c1582; 
    fa fa1582 (s1272, s1273, s1274, s1582, c1582);
    logic s1583 ,c1583; 
    fa fa1583 (c1272, c1273, c1274, s1583, c1583);
    logic s1584 ,c1584; 
    fa fa1584 (s1275, s1276, s1277, s1584, c1584);
    logic s1585 ,c1585; 
    fa fa1585 (c1275, c1276, c1277, s1585, c1585);
    logic s1586 ,c1586; 
    fa fa1586 (s1278, s1279, s1280, s1586, c1586);
    logic s1587 ,c1587; 
    fa fa1587 (c1278, c1279, c1280, s1587, c1587);
    logic s1588 ,c1588; 
    fa fa1588 (s1281, s1282, s1283, s1588, c1588);
    logic s1589 ,c1589; 
    fa fa1589 (c1281, c1282, c1283, s1589, c1589);
    logic s1590 ,c1590; 
    fa fa1590 (s1284, s1285, s1286, s1590, c1590);
    logic s1591 ,c1591; 
    fa fa1591 (c1284, c1285, c1286, s1591, c1591);
    logic s1592 ,c1592; 
    fa fa1592 (s1287, s1288, s1289, s1592, c1592);
    logic s1593 ,c1593; 
    fa fa1593 (c1287, c1288, c1289, s1593, c1593);
    logic s1594 ,c1594; 
    fa fa1594 (s1290, s1291, s1292, s1594, c1594);
    logic s1595 ,c1595; 
    fa fa1595 (c1290, c1291, c1292, s1595, c1595);
    logic s1596 ,c1596; 
    fa fa1596 (s1293, s1294, s1295, s1596, c1596);
    logic s1597 ,c1597; 
    fa fa1597 (c1293, c1294, c1295, s1597, c1597);
    logic s1598 ,c1598; 
    fa fa1598 (s1296, s1297, s1298, s1598, c1598);
    logic s1599 ,c1599; 
    fa fa1599 (c1296, c1297, c1298, s1599, c1599);
    logic s1600 ,c1600; 
    fa fa1600 (s1299, s1300, s1301, s1600, c1600);
    logic s1601 ,c1601; 
    fa fa1601 (c1299, c1300, c1301, s1601, c1601);
    logic s1602 ,c1602; 
    fa fa1602 (s1302, s1303, s1304, s1602, c1602);
    logic s1603 ,c1603; 
    fa fa1603 (c1302, c1303, c1304, s1603, c1603);
    logic s1604 ,c1604; 
    fa fa1604 (s1305, s1306, s1307, s1604, c1604);
    logic s1605 ,c1605; 
    fa fa1605 (c1305, c1306, c1307, s1605, c1605);
    logic s1606 ,c1606; 
    fa fa1606 (s1308, s1309, s1310, s1606, c1606);
    logic s1607 ,c1607; 
    fa fa1607 (c1308, c1309, c1310, s1607, c1607);
    logic s1608 ,c1608; 
    fa fa1608 (s1311, s1312, s1313, s1608, c1608);
    logic s1609 ,c1609; 
    fa fa1609 (c1311, c1312, c1313, s1609, c1609);
    logic s1610 ,c1610; 
    fa fa1610 (s1314, s1315, s1316, s1610, c1610);
    logic s1611 ,c1611; 
    fa fa1611 (c1314, c1315, c1316, s1611, c1611);
    logic s1612 ,c1612; 
    fa fa1612 (s1317, s1318, s1319, s1612, c1612);
    logic s1613 ,c1613; 
    fa fa1613 (c1317, c1318, c1319, s1613, c1613);
    logic s1614 ,c1614; 
    fa fa1614 (s1320, s1321, s1322, s1614, c1614);
    logic s1615 ,c1615; 
    fa fa1615 (c1320, c1321, c1322, s1615, c1615);
    logic s1616 ,c1616; 
    fa fa1616 (s1323, s1324, s1325, s1616, c1616);
    logic s1617 ,c1617; 
    fa fa1617 (c1323, c1324, c1325, s1617, c1617);
    logic s1618 ,c1618; 
    fa fa1618 (s1326, s1327, s1328, s1618, c1618);
    logic s1619 ,c1619; 
    fa fa1619 (c1326, c1327, c1328, s1619, c1619);
    logic s1620 ,c1620; 
    fa fa1620 (s1329, s1330, s1331, s1620, c1620);
    logic s1621 ,c1621; 
    fa fa1621 (c1329, c1330, c1331, s1621, c1621);
    logic s1622 ,c1622; 
    fa fa1622 (s1332, s1333, s1334, s1622, c1622);
    logic s1623 ,c1623; 
    fa fa1623 (c1332, c1333, c1334, s1623, c1623);
    logic s1624 ,c1624; 
    fa fa1624 (s1335, s1336, s1337, s1624, c1624);
    logic s1625 ,c1625; 
    fa fa1625 (c1335, c1336, c1337, s1625, c1625);
    logic s1626 ,c1626; 
    fa fa1626 (s1338, s1339, s1340, s1626, c1626);
    logic s1627 ,c1627; 
    fa fa1627 (c1338, c1339, c1340, s1627, c1627);
    logic s1628 ,c1628; 
    fa fa1628 (s1341, s1342, s1343, s1628, c1628);
    logic s1629 ,c1629; 
    fa fa1629 (c1341, c1342, c1343, s1629, c1629);
    logic s1630 ,c1630; 
    fa fa1630 (s1344, s1345, s1346, s1630, c1630);
    logic s1631 ,c1631; 
    fa fa1631 (c1344, c1345, c1346, s1631, c1631);
    logic s1632 ,c1632; 
    fa fa1632 (s1347, s1348, s1349, s1632, c1632);
    logic s1633 ,c1633; 
    fa fa1633 (c1347, c1348, c1349, s1633, c1633);
    logic s1634 ,c1634; 
    fa fa1634 (s1350, s1351, s1352, s1634, c1634);
    logic s1635 ,c1635; 
    fa fa1635 (c1350, c1351, c1352, s1635, c1635);
    logic s1636 ,c1636; 
    fa fa1636 (s1353, s1354, s1355, s1636, c1636);
    logic s1637 ,c1637; 
    fa fa1637 (c1353, c1354, c1355, s1637, c1637);
    logic s1638 ,c1638; 
    fa fa1638 (s1356, s1357, s1358, s1638, c1638);
    logic s1639 ,c1639; 
    fa fa1639 (c1356, c1357, c1358, s1639, c1639);
    logic s1640 ,c1640; 
    fa fa1640 (s1359, s1360, s1361, s1640, c1640);
    logic s1641 ,c1641; 
    fa fa1641 (c1359, c1360, c1361, s1641, c1641);
    logic s1642 ,c1642; 
    fa fa1642 (s1362, s1363, s1364, s1642, c1642);
    logic s1643 ,c1643; 
    fa fa1643 (c1362, c1363, c1364, s1643, c1643);
    logic s1644 ,c1644; 
    fa fa1644 (s1365, s1366, s1367, s1644, c1644);
    logic s1645 ,c1645; 
    fa fa1645 (c1365, c1366, c1367, s1645, c1645);
    logic s1646 ,c1646; 
    fa fa1646 (s1368, s1369, s1370, s1646, c1646);
    logic s1647 ,c1647; 
    fa fa1647 (c1368, c1369, c1370, s1647, c1647);
    logic s1648 ,c1648; 
    fa fa1648 (s1371, s1372, s1373, s1648, c1648);
    logic s1649 ,c1649; 
    fa fa1649 (c1371, c1372, c1373, s1649, c1649);
    logic s1650 ,c1650; 
    fa fa1650 (s1374, s1375, s1376, s1650, c1650);
    logic s1651 ,c1651; 
    fa fa1651 (c1374, c1375, c1376, s1651, c1651);
    logic s1652 ,c1652; 
    fa fa1652 (s1377, s1378, s1379, s1652, c1652);
    logic s1653 ,c1653; 
    fa fa1653 (c1377, c1378, c1379, s1653, c1653);
    logic s1654 ,c1654; 
    fa fa1654 (s1380, s1381, s1382, s1654, c1654);
    logic s1655 ,c1655; 
    fa fa1655 (c1380, c1381, c1382, s1655, c1655);
    logic s1656 ,c1656; 
    fa fa1656 (s1383, s1384, s1385, s1656, c1656);
    logic s1657 ,c1657; 
    fa fa1657 (c1383, c1384, c1385, s1657, c1657);
    logic s1658 ,c1658; 
    fa fa1658 (s1386, s1387, s1388, s1658, c1658);
    logic s1659 ,c1659; 
    fa fa1659 (c1386, c1387, c1388, s1659, c1659);
    logic s1660 ,c1660; 
    fa fa1660 (s1389, s1390, s1391, s1660, c1660);
    logic s1661 ,c1661; 
    fa fa1661 (c1389, c1390, c1391, s1661, c1661);
    logic s1662 ,c1662; 
    fa fa1662 (s1392, s1393, s1394, s1662, c1662);
    logic s1663 ,c1663; 
    fa fa1663 (c1392, c1393, c1394, s1663, c1663);
    logic s1664 ,c1664; 
    fa fa1664 (s1395, s1396, s1397, s1664, c1664);
    logic s1665 ,c1665; 
    fa fa1665 (c1395, c1396, c1397, s1665, c1665);
    logic s1666 ,c1666; 
    fa fa1666 (s1398, s1399, s1400, s1666, c1666);
    logic s1667 ,c1667; 
    fa fa1667 (c1398, c1399, c1400, s1667, c1667);
    logic s1668 ,c1668; 
    fa fa1668 (s1401, s1402, s1403, s1668, c1668);
    logic s1669 ,c1669; 
    fa fa1669 (c1401, c1402, c1403, s1669, c1669);
    logic s1670 ,c1670; 
    fa fa1670 (s1404, s1405, s1406, s1670, c1670);
    logic s1671 ,c1671; 
    fa fa1671 (c1404, c1405, c1406, s1671, c1671);
    logic s1672 ,c1672; 
    fa fa1672 (s1407, s1408, s1409, s1672, c1672);
    logic s1673 ,c1673; 
    fa fa1673 (c1407, c1408, c1409, s1673, c1673);
    logic s1674 ,c1674; 
    fa fa1674 (s1410, s1411, s1412, s1674, c1674);
    logic s1675 ,c1675; 
    fa fa1675 (c1410, c1411, c1412, s1675, c1675);
    logic s1676 ,c1676; 
    fa fa1676 (s1413, s1414, s1415, s1676, c1676);
    logic s1677 ,c1677; 
    fa fa1677 (c1413, c1414, c1415, s1677, c1677);
    logic s1678 ,c1678; 
    fa fa1678 (s1416, s1417, s1418, s1678, c1678);
    logic s1679 ,c1679; 
    fa fa1679 (c1416, c1417, c1418, s1679, c1679);
    logic s1680 ,c1680; 
    fa fa1680 (s1419, s1420, s1421, s1680, c1680);
    logic s1681 ,c1681; 
    fa fa1681 (c1419, c1420, c1421, s1681, c1681);
    logic s1682 ,c1682; 
    fa fa1682 (s1422, s1423, s1424, s1682, c1682);
    logic s1683 ,c1683; 
    fa fa1683 (c1422, c1423, c1424, s1683, c1683);
    logic s1684 ,c1684; 
    fa fa1684 (s1425, s1426, s1427, s1684, c1684);
    logic s1685 ,c1685; 
    fa fa1685 (c1425, c1426, c1427, s1685, c1685);
    logic s1686 ,c1686; 
    fa fa1686 (s1428, s1429, s1430, s1686, c1686);
    logic s1687 ,c1687; 
    fa fa1687 (c1428, c1429, c1430, s1687, c1687);
    logic s1688 ,c1688; 
    fa fa1688 (s1431, s1432, s1433, s1688, c1688);
    logic s1689 ,c1689; 
    fa fa1689 (c1431, c1432, c1433, s1689, c1689);
    logic s1690 ,c1690; 
    fa fa1690 (s1434, s1435, s1436, s1690, c1690);
    logic s1691 ,c1691; 
    fa fa1691 (c1434, c1435, c1436, s1691, c1691);
    logic s1692 ,c1692; 
    fa fa1692 (s1437, s1438, s1439, s1692, c1692);
    logic s1693 ,c1693; 
    fa fa1693 (c1437, c1438, c1439, s1693, c1693);
    logic s1694 ,c1694; 
    fa fa1694 (s1440, s1441, s1442, s1694, c1694);
    logic s1695 ,c1695; 
    fa fa1695 (c1440, c1441, c1442, s1695, c1695);
    logic s1696 ,c1696; 
    fa fa1696 (s1443, s1444, s1445, s1696, c1696);
    logic s1697 ,c1697; 
    fa fa1697 (c1443, c1444, c1445, s1697, c1697);
    logic s1698 ,c1698; 
    fa fa1698 (s1446, s1447, s1448, s1698, c1698);
    logic s1699 ,c1699; 
    fa fa1699 (c1446, c1447, c1448, s1699, c1699);
    logic s1700 ,c1700; 
    fa fa1700 (s1449, s1450, s1451, s1700, c1700);
    logic s1701 ,c1701; 
    fa fa1701 (c1449, c1450, c1451, s1701, c1701);
    logic s1702 ,c1702; 
    fa fa1702 (s1452, s1453, s1454, s1702, c1702);
    logic s1703 ,c1703; 
    fa fa1703 (c1452, c1453, c1454, s1703, c1703);
    logic s1704 ,c1704; 
    fa fa1704 (s1455, s1456, s1457, s1704, c1704);
    logic s1705 ,c1705; 
    fa fa1705 (c1455, c1456, c1457, s1705, c1705);
    logic s1706 ,c1706; 
    fa fa1706 (s1458, s1459, s1460, s1706, c1706);
    logic s1707 ,c1707; 
    fa fa1707 (c1458, c1459, c1460, s1707, c1707);
    logic s1708 ,c1708; 
    fa fa1708 (s1461, s1462, s1463, s1708, c1708);
    logic s1709 ,c1709; 
    fa fa1709 (c1461, c1462, c1463, s1709, c1709);
    logic s1710 ,c1710; 
    fa fa1710 (s1464, s1465, s1466, s1710, c1710);
    logic s1711 ,c1711; 
    fa fa1711 (c1464, c1465, c1466, s1711, c1711);
    logic s1712 ,c1712; 
    fa fa1712 (s1467, s1468, s1469, s1712, c1712);
    logic s1713 ,c1713; 
    fa fa1713 (c1467, c1468, c1469, s1713, c1713);
    logic s1714 ,c1714; 
    fa fa1714 (s1470, s1471, s1472, s1714, c1714);
    logic s1715 ,c1715; 
    fa fa1715 (c1470, c1471, c1472, s1715, c1715);
    logic s1716 ,c1716; 
    fa fa1716 (s1473, s1474, s1475, s1716, c1716);
    logic s1717 ,c1717; 
    fa fa1717 (c1473, c1474, c1475, s1717, c1717);
    logic s1718 ,c1718; 
    fa fa1718 (s1476, s1477, s1478, s1718, c1718);
    logic s1719 ,c1719; 
    fa fa1719 (c1476, c1477, c1478, s1719, c1719);
    logic s1720 ,c1720; 
    fa fa1720 (s1479, s1480, s1481, s1720, c1720);
    logic s1721 ,c1721; 
    fa fa1721 (c1479, c1480, c1481, s1721, c1721);
    logic s1722 ,c1722; 
    fa fa1722 (s1482, s1483, s1484, s1722, c1722);
    logic s1723 ,c1723; 
    fa fa1723 (c1482, c1483, c1484, s1723, c1723);
    logic s1724 ,c1724; 
    fa fa1724 (s1485, s1486, s1487, s1724, c1724);
    logic s1725 ,c1725; 
    fa fa1725 (c1485, c1486, c1487, s1725, c1725);
    logic s1726 ,c1726; 
    fa fa1726 (s1488, s1489, s1490, s1726, c1726);
    logic s1727 ,c1727; 
    fa fa1727 (c1488, c1489, c1490, s1727, c1727);
    logic s1728 ,c1728; 
    fa fa1728 (s1491, s1492, s1493, s1728, c1728);
    logic s1729 ,c1729; 
    fa fa1729 (c1491, c1492, c1493, s1729, c1729);
    logic s1730 ,c1730; 
    fa fa1730 (s1494, s1495, s1496, s1730, c1730);
    logic s1731 ,c1731; 
    fa fa1731 (c1494, c1495, c1496, s1731, c1731);
    logic s1732 ,c1732; 
    fa fa1732 (s1497, s1498, s1499, s1732, c1732);
    logic s1733 ,c1733; 
    fa fa1733 (c1497, c1498, c1499, s1733, c1733);
    logic s1734 ,c1734; 
    fa fa1734 (s1500, s1501, s1502, s1734, c1734);
    logic s1735 ,c1735; 
    fa fa1735 (c1500, c1501, c1502, s1735, c1735);
    logic s1736 ,c1736; 
    fa fa1736 (s1503, s1504, s1505, s1736, c1736);
    logic s1737 ,c1737; 
    fa fa1737 (c1503, c1504, c1505, s1737, c1737);
    logic s1738 ,c1738; 
    fa fa1738 (s1506, s1507, s1508, s1738, c1738);
    logic s1739 ,c1739; 
    fa fa1739 (c1506, c1507, c1508, s1739, c1739);
    logic s1740 ,c1740; 
    fa fa1740 (s1509, s1510, s1511, s1740, c1740);
    logic s1741 ,c1741; 
    fa fa1741 (c1509, c1510, c1511, s1741, c1741);
    logic s1742 ,c1742; 
    fa fa1742 (s1512, s1513, s1514, s1742, c1742);
    logic s1743 ,c1743; 
    fa fa1743 (c1512, c1513, c1514, s1743, c1743);
    logic s1744 ,c1744; 
    fa fa1744 (s1515, s1516, s1517, s1744, c1744);
    logic s1745 ,c1745; 
    fa fa1745 (c1515, c1516, c1517, s1745, c1745);
    logic s1746 ,c1746; 
    fa fa1746 (s1518, s1519, s1520, s1746, c1746);
    logic s1747 ,c1747; 
    fa fa1747 (c1518, c1519, c1520, s1747, c1747);
    logic s1748 ,c1748; 
    fa fa1748 (s1521, s1522, s1523, s1748, c1748);
    logic s1749 ,c1749; 
    fa fa1749 (c1521, c1522, c1523, s1749, c1749);
    logic s1750 ,c1750; 
    fa fa1750 (s1524, s1525, s1526, s1750, c1750);
    logic s1751 ,c1751; 
    fa fa1751 (c1524, c1525, c1526, s1751, c1751);
    logic s1752 ,c1752; 
    fa fa1752 (s1527, s1528, s1529, s1752, c1752);
    logic s1753 ,c1753; 
    fa fa1753 (c1527, c1528, c1529, s1753, c1753);
    logic s1754 ,c1754; 
    fa fa1754 (s1530, s1531, s1532, s1754, c1754);
    logic s1755 ,c1755; 
    fa fa1755 (pp_31_53, c1530, c1531, s1755, c1755);
    logic s1756 ,c1756; 
    fa fa1756 (c1532, s1533, s1534, s1756, c1756);
    logic s1757 ,c1757; 
    fa fa1757 (pp_30_56, pp_31_54, c1533, s1757, c1757);
    logic s1758 ,c1758; 
    fa fa1758 (c1534, s1535, s1536, s1758, c1758);
    logic s1759 ,c1759; 
    fa fa1759 (pp_29_59, pp_30_57, pp_31_55, s1759, c1759);
    logic s1760 ,c1760; 
    fa fa1760 (c1535, c1536, s1537, s1760, c1760);
    logic s1761 ,c1761; 
    fa fa1761 (pp_28_62, pp_29_60, pp_30_58, s1761, c1761);
    logic s1762 ,c1762; 
    fa fa1762 (pp_31_56, c1537, s1538, s1762, c1762);
    logic s1763 ,c1763; 
    fa fa1763 (pp_27_65, pp_28_63, pp_29_61, s1763, c1763);
    logic s1764 ,c1764; 
    fa fa1764 (pp_30_59, pp_31_57, c1538, s1764, c1764);
    logic s1765 ,c1765; 
    fa fa1765 (const1, pp_28_64, pp_29_62, s1765, c1765);
    logic s1766 ,c1766;
    ha ha1766 (pp_30_60, pp_31_58, s1766, c1766);
    logic s1767 ,c1767; 
    fa fa1767 (pp_28_65, pp_29_63, pp_30_61, s1767, c1767);
    logic s1768 ,c1768;
    ha ha1768 (const1, pp_29_64, s1768, c1768);
    logic s1769 ,c1769;
    ha ha1769 (pp_0_4, pp_1_2, s1769, c1769);
    logic s1770 ,c1770;
    ha ha1770 (pp_0_5, pp_1_3, s1770, c1770);
    logic s1771 ,c1771; 
    fa fa1771 (pp_2_2, pp_3_0, tcomp3, s1771, c1771);
    logic s1772 ,c1772; 
    fa fa1772 (pp_2_3, pp_3_1, c1539, s1772, c1772);
    logic s1773 ,c1773; 
    fa fa1773 (tcomp4, c1540, s1541, s1773, c1773);
    logic s1774 ,c1774; 
    fa fa1774 (c1541, c1542, s1543, s1774, c1774);
    logic s1775 ,c1775; 
    fa fa1775 (c1543, c1544, s1545, s1775, c1775);
    logic s1776 ,c1776; 
    fa fa1776 (c1545, c1546, s1547, s1776, c1776);
    logic s1777 ,c1777; 
    fa fa1777 (c1547, c1548, s1549, s1777, c1777);
    logic s1778 ,c1778; 
    fa fa1778 (c1549, c1550, s1551, s1778, c1778);
    logic s1779 ,c1779; 
    fa fa1779 (c1551, c1552, s1553, s1779, c1779);
    logic s1780 ,c1780; 
    fa fa1780 (c1553, c1554, s1555, s1780, c1780);
    logic s1781 ,c1781; 
    fa fa1781 (c1555, c1556, s1557, s1781, c1781);
    logic s1782 ,c1782; 
    fa fa1782 (c1557, c1558, s1559, s1782, c1782);
    logic s1783 ,c1783; 
    fa fa1783 (c1559, c1560, s1561, s1783, c1783);
    logic s1784 ,c1784; 
    fa fa1784 (c1561, c1562, s1563, s1784, c1784);
    logic s1785 ,c1785; 
    fa fa1785 (c1563, c1564, s1565, s1785, c1785);
    logic s1786 ,c1786; 
    fa fa1786 (c1565, c1566, s1567, s1786, c1786);
    logic s1787 ,c1787; 
    fa fa1787 (c1567, c1568, s1569, s1787, c1787);
    logic s1788 ,c1788; 
    fa fa1788 (c1569, c1570, s1571, s1788, c1788);
    logic s1789 ,c1789; 
    fa fa1789 (c1571, c1572, s1573, s1789, c1789);
    logic s1790 ,c1790; 
    fa fa1790 (c1573, c1574, s1575, s1790, c1790);
    logic s1791 ,c1791; 
    fa fa1791 (c1575, c1576, s1577, s1791, c1791);
    logic s1792 ,c1792; 
    fa fa1792 (c1577, c1578, s1579, s1792, c1792);
    logic s1793 ,c1793; 
    fa fa1793 (c1579, c1580, s1581, s1793, c1793);
    logic s1794 ,c1794; 
    fa fa1794 (c1581, c1582, s1583, s1794, c1794);
    logic s1795 ,c1795; 
    fa fa1795 (c1583, c1584, s1585, s1795, c1795);
    logic s1796 ,c1796; 
    fa fa1796 (c1585, c1586, s1587, s1796, c1796);
    logic s1797 ,c1797; 
    fa fa1797 (c1587, c1588, s1589, s1797, c1797);
    logic s1798 ,c1798; 
    fa fa1798 (c1589, c1590, s1591, s1798, c1798);
    logic s1799 ,c1799; 
    fa fa1799 (c1591, c1592, s1593, s1799, c1799);
    logic s1800 ,c1800; 
    fa fa1800 (c1593, c1594, s1595, s1800, c1800);
    logic s1801 ,c1801; 
    fa fa1801 (c1595, c1596, s1597, s1801, c1801);
    logic s1802 ,c1802; 
    fa fa1802 (c1597, c1598, s1599, s1802, c1802);
    logic s1803 ,c1803; 
    fa fa1803 (c1599, c1600, s1601, s1803, c1803);
    logic s1804 ,c1804; 
    fa fa1804 (c1601, c1602, s1603, s1804, c1804);
    logic s1805 ,c1805; 
    fa fa1805 (c1603, c1604, s1605, s1805, c1805);
    logic s1806 ,c1806; 
    fa fa1806 (c1605, c1606, s1607, s1806, c1806);
    logic s1807 ,c1807; 
    fa fa1807 (c1607, c1608, s1609, s1807, c1807);
    logic s1808 ,c1808; 
    fa fa1808 (c1609, c1610, s1611, s1808, c1808);
    logic s1809 ,c1809; 
    fa fa1809 (c1611, c1612, s1613, s1809, c1809);
    logic s1810 ,c1810; 
    fa fa1810 (c1613, c1614, s1615, s1810, c1810);
    logic s1811 ,c1811; 
    fa fa1811 (c1615, c1616, s1617, s1811, c1811);
    logic s1812 ,c1812; 
    fa fa1812 (c1617, c1618, s1619, s1812, c1812);
    logic s1813 ,c1813; 
    fa fa1813 (c1619, c1620, s1621, s1813, c1813);
    logic s1814 ,c1814; 
    fa fa1814 (c1621, c1622, s1623, s1814, c1814);
    logic s1815 ,c1815; 
    fa fa1815 (c1623, c1624, s1625, s1815, c1815);
    logic s1816 ,c1816; 
    fa fa1816 (c1625, c1626, s1627, s1816, c1816);
    logic s1817 ,c1817; 
    fa fa1817 (c1627, c1628, s1629, s1817, c1817);
    logic s1818 ,c1818; 
    fa fa1818 (c1629, c1630, s1631, s1818, c1818);
    logic s1819 ,c1819; 
    fa fa1819 (c1631, c1632, s1633, s1819, c1819);
    logic s1820 ,c1820; 
    fa fa1820 (c1633, c1634, s1635, s1820, c1820);
    logic s1821 ,c1821; 
    fa fa1821 (c1635, c1636, s1637, s1821, c1821);
    logic s1822 ,c1822; 
    fa fa1822 (c1637, c1638, s1639, s1822, c1822);
    logic s1823 ,c1823; 
    fa fa1823 (c1639, c1640, s1641, s1823, c1823);
    logic s1824 ,c1824; 
    fa fa1824 (c1641, c1642, s1643, s1824, c1824);
    logic s1825 ,c1825; 
    fa fa1825 (c1643, c1644, s1645, s1825, c1825);
    logic s1826 ,c1826; 
    fa fa1826 (c1645, c1646, s1647, s1826, c1826);
    logic s1827 ,c1827; 
    fa fa1827 (c1647, c1648, s1649, s1827, c1827);
    logic s1828 ,c1828; 
    fa fa1828 (c1649, c1650, s1651, s1828, c1828);
    logic s1829 ,c1829; 
    fa fa1829 (c1651, c1652, s1653, s1829, c1829);
    logic s1830 ,c1830; 
    fa fa1830 (c1653, c1654, s1655, s1830, c1830);
    logic s1831 ,c1831; 
    fa fa1831 (c1655, c1656, s1657, s1831, c1831);
    logic s1832 ,c1832; 
    fa fa1832 (c1657, c1658, s1659, s1832, c1832);
    logic s1833 ,c1833; 
    fa fa1833 (c1659, c1660, s1661, s1833, c1833);
    logic s1834 ,c1834; 
    fa fa1834 (c1661, c1662, s1663, s1834, c1834);
    logic s1835 ,c1835; 
    fa fa1835 (c1663, c1664, s1665, s1835, c1835);
    logic s1836 ,c1836; 
    fa fa1836 (c1665, c1666, s1667, s1836, c1836);
    logic s1837 ,c1837; 
    fa fa1837 (c1667, c1668, s1669, s1837, c1837);
    logic s1838 ,c1838; 
    fa fa1838 (c1669, c1670, s1671, s1838, c1838);
    logic s1839 ,c1839; 
    fa fa1839 (c1671, c1672, s1673, s1839, c1839);
    logic s1840 ,c1840; 
    fa fa1840 (c1673, c1674, s1675, s1840, c1840);
    logic s1841 ,c1841; 
    fa fa1841 (c1675, c1676, s1677, s1841, c1841);
    logic s1842 ,c1842; 
    fa fa1842 (c1677, c1678, s1679, s1842, c1842);
    logic s1843 ,c1843; 
    fa fa1843 (c1679, c1680, s1681, s1843, c1843);
    logic s1844 ,c1844; 
    fa fa1844 (c1681, c1682, s1683, s1844, c1844);
    logic s1845 ,c1845; 
    fa fa1845 (c1683, c1684, s1685, s1845, c1845);
    logic s1846 ,c1846; 
    fa fa1846 (c1685, c1686, s1687, s1846, c1846);
    logic s1847 ,c1847; 
    fa fa1847 (c1687, c1688, s1689, s1847, c1847);
    logic s1848 ,c1848; 
    fa fa1848 (c1689, c1690, s1691, s1848, c1848);
    logic s1849 ,c1849; 
    fa fa1849 (c1691, c1692, s1693, s1849, c1849);
    logic s1850 ,c1850; 
    fa fa1850 (c1693, c1694, s1695, s1850, c1850);
    logic s1851 ,c1851; 
    fa fa1851 (c1695, c1696, s1697, s1851, c1851);
    logic s1852 ,c1852; 
    fa fa1852 (c1697, c1698, s1699, s1852, c1852);
    logic s1853 ,c1853; 
    fa fa1853 (c1699, c1700, s1701, s1853, c1853);
    logic s1854 ,c1854; 
    fa fa1854 (c1701, c1702, s1703, s1854, c1854);
    logic s1855 ,c1855; 
    fa fa1855 (c1703, c1704, s1705, s1855, c1855);
    logic s1856 ,c1856; 
    fa fa1856 (c1705, c1706, s1707, s1856, c1856);
    logic s1857 ,c1857; 
    fa fa1857 (c1707, c1708, s1709, s1857, c1857);
    logic s1858 ,c1858; 
    fa fa1858 (c1709, c1710, s1711, s1858, c1858);
    logic s1859 ,c1859; 
    fa fa1859 (c1711, c1712, s1713, s1859, c1859);
    logic s1860 ,c1860; 
    fa fa1860 (c1713, c1714, s1715, s1860, c1860);
    logic s1861 ,c1861; 
    fa fa1861 (c1715, c1716, s1717, s1861, c1861);
    logic s1862 ,c1862; 
    fa fa1862 (c1717, c1718, s1719, s1862, c1862);
    logic s1863 ,c1863; 
    fa fa1863 (c1719, c1720, s1721, s1863, c1863);
    logic s1864 ,c1864; 
    fa fa1864 (c1721, c1722, s1723, s1864, c1864);
    logic s1865 ,c1865; 
    fa fa1865 (c1723, c1724, s1725, s1865, c1865);
    logic s1866 ,c1866; 
    fa fa1866 (c1725, c1726, s1727, s1866, c1866);
    logic s1867 ,c1867; 
    fa fa1867 (c1727, c1728, s1729, s1867, c1867);
    logic s1868 ,c1868; 
    fa fa1868 (c1729, c1730, s1731, s1868, c1868);
    logic s1869 ,c1869; 
    fa fa1869 (c1731, c1732, s1733, s1869, c1869);
    logic s1870 ,c1870; 
    fa fa1870 (c1733, c1734, s1735, s1870, c1870);
    logic s1871 ,c1871; 
    fa fa1871 (c1735, c1736, s1737, s1871, c1871);
    logic s1872 ,c1872; 
    fa fa1872 (c1737, c1738, s1739, s1872, c1872);
    logic s1873 ,c1873; 
    fa fa1873 (c1739, c1740, s1741, s1873, c1873);
    logic s1874 ,c1874; 
    fa fa1874 (c1741, c1742, s1743, s1874, c1874);
    logic s1875 ,c1875; 
    fa fa1875 (c1743, c1744, s1745, s1875, c1875);
    logic s1876 ,c1876; 
    fa fa1876 (c1745, c1746, s1747, s1876, c1876);
    logic s1877 ,c1877; 
    fa fa1877 (c1747, c1748, s1749, s1877, c1877);
    logic s1878 ,c1878; 
    fa fa1878 (c1749, c1750, s1751, s1878, c1878);
    logic s1879 ,c1879; 
    fa fa1879 (c1751, c1752, s1753, s1879, c1879);
    logic s1880 ,c1880; 
    fa fa1880 (c1753, c1754, s1755, s1880, c1880);
    logic s1881 ,c1881; 
    fa fa1881 (c1755, c1756, s1757, s1881, c1881);
    logic s1882 ,c1882; 
    fa fa1882 (c1757, c1758, s1759, s1882, c1882);
    logic s1883 ,c1883; 
    fa fa1883 (c1759, c1760, s1761, s1883, c1883);
    logic s1884 ,c1884; 
    fa fa1884 (c1761, c1762, s1763, s1884, c1884);
    logic s1885 ,c1885; 
    fa fa1885 (c1763, c1764, s1765, s1885, c1885);
    logic s1886 ,c1886; 
    fa fa1886 (pp_31_59, c1765, c1766, s1886, c1886);
    logic s1887 ,c1887; 
    fa fa1887 (pp_30_62, pp_31_60, c1767, s1887, c1887);
    logic s1888 ,c1888; 
    fa fa1888 (pp_29_65, pp_30_63, pp_31_61, s1888, c1888);
    logic s1889 ,c1889;
    ha ha1889 (const1, pp_30_64, s1889, c1889);
    logic s1890 ,c1890;
    ha ha1890 (pp_0_2, pp_1_0, s1890, c1890);
    logic s1891 ,c1891;
    ha ha1891 (pp_0_3, pp_1_1, s1891, c1891);
    logic s1892 ,c1892; 
    fa fa1892 (pp_2_0, tcomp2, s1769, s1892, c1892);
    logic s1893 ,c1893; 
    fa fa1893 (pp_2_1, c1769, s1770, s1893, c1893);
    logic s1894 ,c1894; 
    fa fa1894 (s1539, c1770, s1771, s1894, c1894);
    logic s1895 ,c1895; 
    fa fa1895 (s1540, c1771, s1772, s1895, c1895);
    logic s1896 ,c1896; 
    fa fa1896 (s1542, c1772, s1773, s1896, c1896);
    logic s1897 ,c1897; 
    fa fa1897 (s1544, c1773, s1774, s1897, c1897);
    logic s1898 ,c1898; 
    fa fa1898 (s1546, c1774, s1775, s1898, c1898);
    logic s1899 ,c1899; 
    fa fa1899 (s1548, c1775, s1776, s1899, c1899);
    logic s1900 ,c1900; 
    fa fa1900 (s1550, c1776, s1777, s1900, c1900);
    logic s1901 ,c1901; 
    fa fa1901 (s1552, c1777, s1778, s1901, c1901);
    logic s1902 ,c1902; 
    fa fa1902 (s1554, c1778, s1779, s1902, c1902);
    logic s1903 ,c1903; 
    fa fa1903 (s1556, c1779, s1780, s1903, c1903);
    logic s1904 ,c1904; 
    fa fa1904 (s1558, c1780, s1781, s1904, c1904);
    logic s1905 ,c1905; 
    fa fa1905 (s1560, c1781, s1782, s1905, c1905);
    logic s1906 ,c1906; 
    fa fa1906 (s1562, c1782, s1783, s1906, c1906);
    logic s1907 ,c1907; 
    fa fa1907 (s1564, c1783, s1784, s1907, c1907);
    logic s1908 ,c1908; 
    fa fa1908 (s1566, c1784, s1785, s1908, c1908);
    logic s1909 ,c1909; 
    fa fa1909 (s1568, c1785, s1786, s1909, c1909);
    logic s1910 ,c1910; 
    fa fa1910 (s1570, c1786, s1787, s1910, c1910);
    logic s1911 ,c1911; 
    fa fa1911 (s1572, c1787, s1788, s1911, c1911);
    logic s1912 ,c1912; 
    fa fa1912 (s1574, c1788, s1789, s1912, c1912);
    logic s1913 ,c1913; 
    fa fa1913 (s1576, c1789, s1790, s1913, c1913);
    logic s1914 ,c1914; 
    fa fa1914 (s1578, c1790, s1791, s1914, c1914);
    logic s1915 ,c1915; 
    fa fa1915 (s1580, c1791, s1792, s1915, c1915);
    logic s1916 ,c1916; 
    fa fa1916 (s1582, c1792, s1793, s1916, c1916);
    logic s1917 ,c1917; 
    fa fa1917 (s1584, c1793, s1794, s1917, c1917);
    logic s1918 ,c1918; 
    fa fa1918 (s1586, c1794, s1795, s1918, c1918);
    logic s1919 ,c1919; 
    fa fa1919 (s1588, c1795, s1796, s1919, c1919);
    logic s1920 ,c1920; 
    fa fa1920 (s1590, c1796, s1797, s1920, c1920);
    logic s1921 ,c1921; 
    fa fa1921 (s1592, c1797, s1798, s1921, c1921);
    logic s1922 ,c1922; 
    fa fa1922 (s1594, c1798, s1799, s1922, c1922);
    logic s1923 ,c1923; 
    fa fa1923 (s1596, c1799, s1800, s1923, c1923);
    logic s1924 ,c1924; 
    fa fa1924 (s1598, c1800, s1801, s1924, c1924);
    logic s1925 ,c1925; 
    fa fa1925 (s1600, c1801, s1802, s1925, c1925);
    logic s1926 ,c1926; 
    fa fa1926 (s1602, c1802, s1803, s1926, c1926);
    logic s1927 ,c1927; 
    fa fa1927 (s1604, c1803, s1804, s1927, c1927);
    logic s1928 ,c1928; 
    fa fa1928 (s1606, c1804, s1805, s1928, c1928);
    logic s1929 ,c1929; 
    fa fa1929 (s1608, c1805, s1806, s1929, c1929);
    logic s1930 ,c1930; 
    fa fa1930 (s1610, c1806, s1807, s1930, c1930);
    logic s1931 ,c1931; 
    fa fa1931 (s1612, c1807, s1808, s1931, c1931);
    logic s1932 ,c1932; 
    fa fa1932 (s1614, c1808, s1809, s1932, c1932);
    logic s1933 ,c1933; 
    fa fa1933 (s1616, c1809, s1810, s1933, c1933);
    logic s1934 ,c1934; 
    fa fa1934 (s1618, c1810, s1811, s1934, c1934);
    logic s1935 ,c1935; 
    fa fa1935 (s1620, c1811, s1812, s1935, c1935);
    logic s1936 ,c1936; 
    fa fa1936 (s1622, c1812, s1813, s1936, c1936);
    logic s1937 ,c1937; 
    fa fa1937 (s1624, c1813, s1814, s1937, c1937);
    logic s1938 ,c1938; 
    fa fa1938 (s1626, c1814, s1815, s1938, c1938);
    logic s1939 ,c1939; 
    fa fa1939 (s1628, c1815, s1816, s1939, c1939);
    logic s1940 ,c1940; 
    fa fa1940 (s1630, c1816, s1817, s1940, c1940);
    logic s1941 ,c1941; 
    fa fa1941 (s1632, c1817, s1818, s1941, c1941);
    logic s1942 ,c1942; 
    fa fa1942 (s1634, c1818, s1819, s1942, c1942);
    logic s1943 ,c1943; 
    fa fa1943 (s1636, c1819, s1820, s1943, c1943);
    logic s1944 ,c1944; 
    fa fa1944 (s1638, c1820, s1821, s1944, c1944);
    logic s1945 ,c1945; 
    fa fa1945 (s1640, c1821, s1822, s1945, c1945);
    logic s1946 ,c1946; 
    fa fa1946 (s1642, c1822, s1823, s1946, c1946);
    logic s1947 ,c1947; 
    fa fa1947 (s1644, c1823, s1824, s1947, c1947);
    logic s1948 ,c1948; 
    fa fa1948 (s1646, c1824, s1825, s1948, c1948);
    logic s1949 ,c1949; 
    fa fa1949 (s1648, c1825, s1826, s1949, c1949);
    logic s1950 ,c1950; 
    fa fa1950 (s1650, c1826, s1827, s1950, c1950);
    logic s1951 ,c1951; 
    fa fa1951 (s1652, c1827, s1828, s1951, c1951);
    logic s1952 ,c1952; 
    fa fa1952 (s1654, c1828, s1829, s1952, c1952);
    logic s1953 ,c1953; 
    fa fa1953 (s1656, c1829, s1830, s1953, c1953);
    logic s1954 ,c1954; 
    fa fa1954 (s1658, c1830, s1831, s1954, c1954);
    logic s1955 ,c1955; 
    fa fa1955 (s1660, c1831, s1832, s1955, c1955);
    logic s1956 ,c1956; 
    fa fa1956 (s1662, c1832, s1833, s1956, c1956);
    logic s1957 ,c1957; 
    fa fa1957 (s1664, c1833, s1834, s1957, c1957);
    logic s1958 ,c1958; 
    fa fa1958 (s1666, c1834, s1835, s1958, c1958);
    logic s1959 ,c1959; 
    fa fa1959 (s1668, c1835, s1836, s1959, c1959);
    logic s1960 ,c1960; 
    fa fa1960 (s1670, c1836, s1837, s1960, c1960);
    logic s1961 ,c1961; 
    fa fa1961 (s1672, c1837, s1838, s1961, c1961);
    logic s1962 ,c1962; 
    fa fa1962 (s1674, c1838, s1839, s1962, c1962);
    logic s1963 ,c1963; 
    fa fa1963 (s1676, c1839, s1840, s1963, c1963);
    logic s1964 ,c1964; 
    fa fa1964 (s1678, c1840, s1841, s1964, c1964);
    logic s1965 ,c1965; 
    fa fa1965 (s1680, c1841, s1842, s1965, c1965);
    logic s1966 ,c1966; 
    fa fa1966 (s1682, c1842, s1843, s1966, c1966);
    logic s1967 ,c1967; 
    fa fa1967 (s1684, c1843, s1844, s1967, c1967);
    logic s1968 ,c1968; 
    fa fa1968 (s1686, c1844, s1845, s1968, c1968);
    logic s1969 ,c1969; 
    fa fa1969 (s1688, c1845, s1846, s1969, c1969);
    logic s1970 ,c1970; 
    fa fa1970 (s1690, c1846, s1847, s1970, c1970);
    logic s1971 ,c1971; 
    fa fa1971 (s1692, c1847, s1848, s1971, c1971);
    logic s1972 ,c1972; 
    fa fa1972 (s1694, c1848, s1849, s1972, c1972);
    logic s1973 ,c1973; 
    fa fa1973 (s1696, c1849, s1850, s1973, c1973);
    logic s1974 ,c1974; 
    fa fa1974 (s1698, c1850, s1851, s1974, c1974);
    logic s1975 ,c1975; 
    fa fa1975 (s1700, c1851, s1852, s1975, c1975);
    logic s1976 ,c1976; 
    fa fa1976 (s1702, c1852, s1853, s1976, c1976);
    logic s1977 ,c1977; 
    fa fa1977 (s1704, c1853, s1854, s1977, c1977);
    logic s1978 ,c1978; 
    fa fa1978 (s1706, c1854, s1855, s1978, c1978);
    logic s1979 ,c1979; 
    fa fa1979 (s1708, c1855, s1856, s1979, c1979);
    logic s1980 ,c1980; 
    fa fa1980 (s1710, c1856, s1857, s1980, c1980);
    logic s1981 ,c1981; 
    fa fa1981 (s1712, c1857, s1858, s1981, c1981);
    logic s1982 ,c1982; 
    fa fa1982 (s1714, c1858, s1859, s1982, c1982);
    logic s1983 ,c1983; 
    fa fa1983 (s1716, c1859, s1860, s1983, c1983);
    logic s1984 ,c1984; 
    fa fa1984 (s1718, c1860, s1861, s1984, c1984);
    logic s1985 ,c1985; 
    fa fa1985 (s1720, c1861, s1862, s1985, c1985);
    logic s1986 ,c1986; 
    fa fa1986 (s1722, c1862, s1863, s1986, c1986);
    logic s1987 ,c1987; 
    fa fa1987 (s1724, c1863, s1864, s1987, c1987);
    logic s1988 ,c1988; 
    fa fa1988 (s1726, c1864, s1865, s1988, c1988);
    logic s1989 ,c1989; 
    fa fa1989 (s1728, c1865, s1866, s1989, c1989);
    logic s1990 ,c1990; 
    fa fa1990 (s1730, c1866, s1867, s1990, c1990);
    logic s1991 ,c1991; 
    fa fa1991 (s1732, c1867, s1868, s1991, c1991);
    logic s1992 ,c1992; 
    fa fa1992 (s1734, c1868, s1869, s1992, c1992);
    logic s1993 ,c1993; 
    fa fa1993 (s1736, c1869, s1870, s1993, c1993);
    logic s1994 ,c1994; 
    fa fa1994 (s1738, c1870, s1871, s1994, c1994);
    logic s1995 ,c1995; 
    fa fa1995 (s1740, c1871, s1872, s1995, c1995);
    logic s1996 ,c1996; 
    fa fa1996 (s1742, c1872, s1873, s1996, c1996);
    logic s1997 ,c1997; 
    fa fa1997 (s1744, c1873, s1874, s1997, c1997);
    logic s1998 ,c1998; 
    fa fa1998 (s1746, c1874, s1875, s1998, c1998);
    logic s1999 ,c1999; 
    fa fa1999 (s1748, c1875, s1876, s1999, c1999);
    logic s2000 ,c2000; 
    fa fa2000 (s1750, c1876, s1877, s2000, c2000);
    logic s2001 ,c2001; 
    fa fa2001 (s1752, c1877, s1878, s2001, c2001);
    logic s2002 ,c2002; 
    fa fa2002 (s1754, c1878, s1879, s2002, c2002);
    logic s2003 ,c2003; 
    fa fa2003 (s1756, c1879, s1880, s2003, c2003);
    logic s2004 ,c2004; 
    fa fa2004 (s1758, c1880, s1881, s2004, c2004);
    logic s2005 ,c2005; 
    fa fa2005 (s1760, c1881, s1882, s2005, c2005);
    logic s2006 ,c2006; 
    fa fa2006 (s1762, c1882, s1883, s2006, c2006);
    logic s2007 ,c2007; 
    fa fa2007 (s1764, c1883, s1884, s2007, c2007);
    logic s2008 ,c2008; 
    fa fa2008 (s1766, c1884, s1885, s2008, c2008);
    logic s2009 ,c2009; 
    fa fa2009 (s1767, c1885, s1886, s2009, c2009);
    logic s2010 ,c2010; 
    fa fa2010 (s1768, c1886, s1887, s2010, c2010);
    logic s2011 ,c2011; 
    fa fa2011 (c1768, c1887, s1888, s2011, c2011);
    logic s2012 ,c2012; 
    fa fa2012 (pp_31_62, c1888, s1889, s2012, c2012);
    logic s2013 ,c2013; 
    fa fa2013 (pp_30_65, pp_31_63, c1889, s2013, c2013);
    logic s2014 ,c2014;
    ha ha2014 (const1, pp_31_64, s2014, c2014);
    logic [128:0] adder_result;
    HC_128 final_adder ({pp_31_65, c2013, c2012, c2011, c2010, c2009, c2008, c2007, c2006, c2005, c2004, c2003, c2002, c2001, c2000, c1999, c1998, c1997, c1996, c1995, c1994, c1993, c1992, c1991, c1990, c1989, c1988, c1987, c1986, c1985, c1984, c1983, c1982, c1981, c1980, c1979, c1978, c1977, c1976, c1975, c1974, c1973, c1972, c1971, c1970, c1969, c1968, c1967, c1966, c1965, c1964, c1963, c1962, c1961, c1960, c1959, c1958, c1957, c1956, c1955, c1954, c1953, c1952, c1951, c1950, c1949, c1948, c1947, c1946, c1945, c1944, c1943, c1942, c1941, c1940, c1939, c1938, c1937, c1936, c1935, c1934, c1933, c1932, c1931, c1930, c1929, c1928, c1927, c1926, c1925, c1924, c1923, c1922, c1921, c1920, c1919, c1918, c1917, c1916, c1915, c1914, c1913, c1912, c1911, c1910, c1909, c1908, c1907, c1906, c1905, c1904, c1903, c1902, c1901, c1900, c1899, c1898, c1897, c1896, c1895, c1894, c1893, c1892, c1891, c1890, tcomp1, pp_0_1, pp_0_0 }, {c2014, s2014, s2013, s2012, s2011, s2010, s2009, s2008, s2007, s2006, s2005, s2004, s2003, s2002, s2001, s2000, s1999, s1998, s1997, s1996, s1995, s1994, s1993, s1992, s1991, s1990, s1989, s1988, s1987, s1986, s1985, s1984, s1983, s1982, s1981, s1980, s1979, s1978, s1977, s1976, s1975, s1974, s1973, s1972, s1971, s1970, s1969, s1968, s1967, s1966, s1965, s1964, s1963, s1962, s1961, s1960, s1959, s1958, s1957, s1956, s1955, s1954, s1953, s1952, s1951, s1950, s1949, s1948, s1947, s1946, s1945, s1944, s1943, s1942, s1941, s1940, s1939, s1938, s1937, s1936, s1935, s1934, s1933, s1932, s1931, s1930, s1929, s1928, s1927, s1926, s1925, s1924, s1923, s1922, s1921, s1920, s1919, s1918, s1917, s1916, s1915, s1914, s1913, s1912, s1911, s1910, s1909, s1908, s1907, s1906, s1905, s1904, s1903, s1902, s1901, s1900, s1899, s1898, s1897, s1896, s1895, s1894, s1893, s1892, s1891, s1890, 1'b0, tcomp0 }, adder_result );
    assign result[127:0] = adder_result[127:0];
    endmodule



module HC_128 ( 
        input logic [127:0] IN1,
        input logic [127:0] IN2,
        output logic [128:0] OUT);
    
    wire logic [127:0] p_0;
    wire logic [127:0] g_0;
    assign g_0 = IN1 & IN2;
    assign p_0 = IN1 ^ IN2;
    
    // HC stage 1
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_3;
    wire logic g_1_3;
    assign p_1_3 = p_0[3] & p_0[2];
    assign g_1_3 = (p_0[3] & g_0[2]) | g_0[3];
    wire logic p_1_5;
    wire logic g_1_5;
    assign p_1_5 = p_0[5] & p_0[4];
    assign g_1_5 = (p_0[5] & g_0[4]) | g_0[5];
    wire logic p_1_7;
    wire logic g_1_7;
    assign p_1_7 = p_0[7] & p_0[6];
    assign g_1_7 = (p_0[7] & g_0[6]) | g_0[7];
    wire logic p_1_9;
    wire logic g_1_9;
    assign p_1_9 = p_0[9] & p_0[8];
    assign g_1_9 = (p_0[9] & g_0[8]) | g_0[9];
    wire logic p_1_11;
    wire logic g_1_11;
    assign p_1_11 = p_0[11] & p_0[10];
    assign g_1_11 = (p_0[11] & g_0[10]) | g_0[11];
    wire logic p_1_13;
    wire logic g_1_13;
    assign p_1_13 = p_0[13] & p_0[12];
    assign g_1_13 = (p_0[13] & g_0[12]) | g_0[13];
    wire logic p_1_15;
    wire logic g_1_15;
    assign p_1_15 = p_0[15] & p_0[14];
    assign g_1_15 = (p_0[15] & g_0[14]) | g_0[15];
    wire logic p_1_17;
    wire logic g_1_17;
    assign p_1_17 = p_0[17] & p_0[16];
    assign g_1_17 = (p_0[17] & g_0[16]) | g_0[17];
    wire logic p_1_19;
    wire logic g_1_19;
    assign p_1_19 = p_0[19] & p_0[18];
    assign g_1_19 = (p_0[19] & g_0[18]) | g_0[19];
    wire logic p_1_21;
    wire logic g_1_21;
    assign p_1_21 = p_0[21] & p_0[20];
    assign g_1_21 = (p_0[21] & g_0[20]) | g_0[21];
    wire logic p_1_23;
    wire logic g_1_23;
    assign p_1_23 = p_0[23] & p_0[22];
    assign g_1_23 = (p_0[23] & g_0[22]) | g_0[23];
    wire logic p_1_25;
    wire logic g_1_25;
    assign p_1_25 = p_0[25] & p_0[24];
    assign g_1_25 = (p_0[25] & g_0[24]) | g_0[25];
    wire logic p_1_27;
    wire logic g_1_27;
    assign p_1_27 = p_0[27] & p_0[26];
    assign g_1_27 = (p_0[27] & g_0[26]) | g_0[27];
    wire logic p_1_29;
    wire logic g_1_29;
    assign p_1_29 = p_0[29] & p_0[28];
    assign g_1_29 = (p_0[29] & g_0[28]) | g_0[29];
    wire logic p_1_31;
    wire logic g_1_31;
    assign p_1_31 = p_0[31] & p_0[30];
    assign g_1_31 = (p_0[31] & g_0[30]) | g_0[31];
    wire logic p_1_33;
    wire logic g_1_33;
    assign p_1_33 = p_0[33] & p_0[32];
    assign g_1_33 = (p_0[33] & g_0[32]) | g_0[33];
    wire logic p_1_35;
    wire logic g_1_35;
    assign p_1_35 = p_0[35] & p_0[34];
    assign g_1_35 = (p_0[35] & g_0[34]) | g_0[35];
    wire logic p_1_37;
    wire logic g_1_37;
    assign p_1_37 = p_0[37] & p_0[36];
    assign g_1_37 = (p_0[37] & g_0[36]) | g_0[37];
    wire logic p_1_39;
    wire logic g_1_39;
    assign p_1_39 = p_0[39] & p_0[38];
    assign g_1_39 = (p_0[39] & g_0[38]) | g_0[39];
    wire logic p_1_41;
    wire logic g_1_41;
    assign p_1_41 = p_0[41] & p_0[40];
    assign g_1_41 = (p_0[41] & g_0[40]) | g_0[41];
    wire logic p_1_43;
    wire logic g_1_43;
    assign p_1_43 = p_0[43] & p_0[42];
    assign g_1_43 = (p_0[43] & g_0[42]) | g_0[43];
    wire logic p_1_45;
    wire logic g_1_45;
    assign p_1_45 = p_0[45] & p_0[44];
    assign g_1_45 = (p_0[45] & g_0[44]) | g_0[45];
    wire logic p_1_47;
    wire logic g_1_47;
    assign p_1_47 = p_0[47] & p_0[46];
    assign g_1_47 = (p_0[47] & g_0[46]) | g_0[47];
    wire logic p_1_49;
    wire logic g_1_49;
    assign p_1_49 = p_0[49] & p_0[48];
    assign g_1_49 = (p_0[49] & g_0[48]) | g_0[49];
    wire logic p_1_51;
    wire logic g_1_51;
    assign p_1_51 = p_0[51] & p_0[50];
    assign g_1_51 = (p_0[51] & g_0[50]) | g_0[51];
    wire logic p_1_53;
    wire logic g_1_53;
    assign p_1_53 = p_0[53] & p_0[52];
    assign g_1_53 = (p_0[53] & g_0[52]) | g_0[53];
    wire logic p_1_55;
    wire logic g_1_55;
    assign p_1_55 = p_0[55] & p_0[54];
    assign g_1_55 = (p_0[55] & g_0[54]) | g_0[55];
    wire logic p_1_57;
    wire logic g_1_57;
    assign p_1_57 = p_0[57] & p_0[56];
    assign g_1_57 = (p_0[57] & g_0[56]) | g_0[57];
    wire logic p_1_59;
    wire logic g_1_59;
    assign p_1_59 = p_0[59] & p_0[58];
    assign g_1_59 = (p_0[59] & g_0[58]) | g_0[59];
    wire logic p_1_61;
    wire logic g_1_61;
    assign p_1_61 = p_0[61] & p_0[60];
    assign g_1_61 = (p_0[61] & g_0[60]) | g_0[61];
    wire logic p_1_63;
    wire logic g_1_63;
    assign p_1_63 = p_0[63] & p_0[62];
    assign g_1_63 = (p_0[63] & g_0[62]) | g_0[63];
    wire logic p_1_65;
    wire logic g_1_65;
    assign p_1_65 = p_0[65] & p_0[64];
    assign g_1_65 = (p_0[65] & g_0[64]) | g_0[65];
    wire logic p_1_67;
    wire logic g_1_67;
    assign p_1_67 = p_0[67] & p_0[66];
    assign g_1_67 = (p_0[67] & g_0[66]) | g_0[67];
    wire logic p_1_69;
    wire logic g_1_69;
    assign p_1_69 = p_0[69] & p_0[68];
    assign g_1_69 = (p_0[69] & g_0[68]) | g_0[69];
    wire logic p_1_71;
    wire logic g_1_71;
    assign p_1_71 = p_0[71] & p_0[70];
    assign g_1_71 = (p_0[71] & g_0[70]) | g_0[71];
    wire logic p_1_73;
    wire logic g_1_73;
    assign p_1_73 = p_0[73] & p_0[72];
    assign g_1_73 = (p_0[73] & g_0[72]) | g_0[73];
    wire logic p_1_75;
    wire logic g_1_75;
    assign p_1_75 = p_0[75] & p_0[74];
    assign g_1_75 = (p_0[75] & g_0[74]) | g_0[75];
    wire logic p_1_77;
    wire logic g_1_77;
    assign p_1_77 = p_0[77] & p_0[76];
    assign g_1_77 = (p_0[77] & g_0[76]) | g_0[77];
    wire logic p_1_79;
    wire logic g_1_79;
    assign p_1_79 = p_0[79] & p_0[78];
    assign g_1_79 = (p_0[79] & g_0[78]) | g_0[79];
    wire logic p_1_81;
    wire logic g_1_81;
    assign p_1_81 = p_0[81] & p_0[80];
    assign g_1_81 = (p_0[81] & g_0[80]) | g_0[81];
    wire logic p_1_83;
    wire logic g_1_83;
    assign p_1_83 = p_0[83] & p_0[82];
    assign g_1_83 = (p_0[83] & g_0[82]) | g_0[83];
    wire logic p_1_85;
    wire logic g_1_85;
    assign p_1_85 = p_0[85] & p_0[84];
    assign g_1_85 = (p_0[85] & g_0[84]) | g_0[85];
    wire logic p_1_87;
    wire logic g_1_87;
    assign p_1_87 = p_0[87] & p_0[86];
    assign g_1_87 = (p_0[87] & g_0[86]) | g_0[87];
    wire logic p_1_89;
    wire logic g_1_89;
    assign p_1_89 = p_0[89] & p_0[88];
    assign g_1_89 = (p_0[89] & g_0[88]) | g_0[89];
    wire logic p_1_91;
    wire logic g_1_91;
    assign p_1_91 = p_0[91] & p_0[90];
    assign g_1_91 = (p_0[91] & g_0[90]) | g_0[91];
    wire logic p_1_93;
    wire logic g_1_93;
    assign p_1_93 = p_0[93] & p_0[92];
    assign g_1_93 = (p_0[93] & g_0[92]) | g_0[93];
    wire logic p_1_95;
    wire logic g_1_95;
    assign p_1_95 = p_0[95] & p_0[94];
    assign g_1_95 = (p_0[95] & g_0[94]) | g_0[95];
    wire logic p_1_97;
    wire logic g_1_97;
    assign p_1_97 = p_0[97] & p_0[96];
    assign g_1_97 = (p_0[97] & g_0[96]) | g_0[97];
    wire logic p_1_99;
    wire logic g_1_99;
    assign p_1_99 = p_0[99] & p_0[98];
    assign g_1_99 = (p_0[99] & g_0[98]) | g_0[99];
    wire logic p_1_101;
    wire logic g_1_101;
    assign p_1_101 = p_0[101] & p_0[100];
    assign g_1_101 = (p_0[101] & g_0[100]) | g_0[101];
    wire logic p_1_103;
    wire logic g_1_103;
    assign p_1_103 = p_0[103] & p_0[102];
    assign g_1_103 = (p_0[103] & g_0[102]) | g_0[103];
    wire logic p_1_105;
    wire logic g_1_105;
    assign p_1_105 = p_0[105] & p_0[104];
    assign g_1_105 = (p_0[105] & g_0[104]) | g_0[105];
    wire logic p_1_107;
    wire logic g_1_107;
    assign p_1_107 = p_0[107] & p_0[106];
    assign g_1_107 = (p_0[107] & g_0[106]) | g_0[107];
    wire logic p_1_109;
    wire logic g_1_109;
    assign p_1_109 = p_0[109] & p_0[108];
    assign g_1_109 = (p_0[109] & g_0[108]) | g_0[109];
    wire logic p_1_111;
    wire logic g_1_111;
    assign p_1_111 = p_0[111] & p_0[110];
    assign g_1_111 = (p_0[111] & g_0[110]) | g_0[111];
    wire logic p_1_113;
    wire logic g_1_113;
    assign p_1_113 = p_0[113] & p_0[112];
    assign g_1_113 = (p_0[113] & g_0[112]) | g_0[113];
    wire logic p_1_115;
    wire logic g_1_115;
    assign p_1_115 = p_0[115] & p_0[114];
    assign g_1_115 = (p_0[115] & g_0[114]) | g_0[115];
    wire logic p_1_117;
    wire logic g_1_117;
    assign p_1_117 = p_0[117] & p_0[116];
    assign g_1_117 = (p_0[117] & g_0[116]) | g_0[117];
    wire logic p_1_119;
    wire logic g_1_119;
    assign p_1_119 = p_0[119] & p_0[118];
    assign g_1_119 = (p_0[119] & g_0[118]) | g_0[119];
    wire logic p_1_121;
    wire logic g_1_121;
    assign p_1_121 = p_0[121] & p_0[120];
    assign g_1_121 = (p_0[121] & g_0[120]) | g_0[121];
    wire logic p_1_123;
    wire logic g_1_123;
    assign p_1_123 = p_0[123] & p_0[122];
    assign g_1_123 = (p_0[123] & g_0[122]) | g_0[123];
    wire logic p_1_125;
    wire logic g_1_125;
    assign p_1_125 = p_0[125] & p_0[124];
    assign g_1_125 = (p_0[125] & g_0[124]) | g_0[125];
    wire logic p_1_127;
    wire logic g_1_127;
    assign p_1_127 = p_0[127] & p_0[126];
    assign g_1_127 = (p_0[127] & g_0[126]) | g_0[127];
    
    // HC stage 2
    wire logic p_2_3;
    wire logic g_2_3;
    assign p_2_3 = p_1_3 & p_1_1;
    assign g_2_3 = (p_1_3 & g_1_1) | g_1_3;
    wire logic p_2_5;
    wire logic g_2_5;
    assign p_2_5 = p_1_5 & p_1_3;
    assign g_2_5 = (p_1_5 & g_1_3) | g_1_5;
    wire logic p_2_7;
    wire logic g_2_7;
    assign p_2_7 = p_1_7 & p_1_5;
    assign g_2_7 = (p_1_7 & g_1_5) | g_1_7;
    wire logic p_2_9;
    wire logic g_2_9;
    assign p_2_9 = p_1_9 & p_1_7;
    assign g_2_9 = (p_1_9 & g_1_7) | g_1_9;
    wire logic p_2_11;
    wire logic g_2_11;
    assign p_2_11 = p_1_11 & p_1_9;
    assign g_2_11 = (p_1_11 & g_1_9) | g_1_11;
    wire logic p_2_13;
    wire logic g_2_13;
    assign p_2_13 = p_1_13 & p_1_11;
    assign g_2_13 = (p_1_13 & g_1_11) | g_1_13;
    wire logic p_2_15;
    wire logic g_2_15;
    assign p_2_15 = p_1_15 & p_1_13;
    assign g_2_15 = (p_1_15 & g_1_13) | g_1_15;
    wire logic p_2_17;
    wire logic g_2_17;
    assign p_2_17 = p_1_17 & p_1_15;
    assign g_2_17 = (p_1_17 & g_1_15) | g_1_17;
    wire logic p_2_19;
    wire logic g_2_19;
    assign p_2_19 = p_1_19 & p_1_17;
    assign g_2_19 = (p_1_19 & g_1_17) | g_1_19;
    wire logic p_2_21;
    wire logic g_2_21;
    assign p_2_21 = p_1_21 & p_1_19;
    assign g_2_21 = (p_1_21 & g_1_19) | g_1_21;
    wire logic p_2_23;
    wire logic g_2_23;
    assign p_2_23 = p_1_23 & p_1_21;
    assign g_2_23 = (p_1_23 & g_1_21) | g_1_23;
    wire logic p_2_25;
    wire logic g_2_25;
    assign p_2_25 = p_1_25 & p_1_23;
    assign g_2_25 = (p_1_25 & g_1_23) | g_1_25;
    wire logic p_2_27;
    wire logic g_2_27;
    assign p_2_27 = p_1_27 & p_1_25;
    assign g_2_27 = (p_1_27 & g_1_25) | g_1_27;
    wire logic p_2_29;
    wire logic g_2_29;
    assign p_2_29 = p_1_29 & p_1_27;
    assign g_2_29 = (p_1_29 & g_1_27) | g_1_29;
    wire logic p_2_31;
    wire logic g_2_31;
    assign p_2_31 = p_1_31 & p_1_29;
    assign g_2_31 = (p_1_31 & g_1_29) | g_1_31;
    wire logic p_2_33;
    wire logic g_2_33;
    assign p_2_33 = p_1_33 & p_1_31;
    assign g_2_33 = (p_1_33 & g_1_31) | g_1_33;
    wire logic p_2_35;
    wire logic g_2_35;
    assign p_2_35 = p_1_35 & p_1_33;
    assign g_2_35 = (p_1_35 & g_1_33) | g_1_35;
    wire logic p_2_37;
    wire logic g_2_37;
    assign p_2_37 = p_1_37 & p_1_35;
    assign g_2_37 = (p_1_37 & g_1_35) | g_1_37;
    wire logic p_2_39;
    wire logic g_2_39;
    assign p_2_39 = p_1_39 & p_1_37;
    assign g_2_39 = (p_1_39 & g_1_37) | g_1_39;
    wire logic p_2_41;
    wire logic g_2_41;
    assign p_2_41 = p_1_41 & p_1_39;
    assign g_2_41 = (p_1_41 & g_1_39) | g_1_41;
    wire logic p_2_43;
    wire logic g_2_43;
    assign p_2_43 = p_1_43 & p_1_41;
    assign g_2_43 = (p_1_43 & g_1_41) | g_1_43;
    wire logic p_2_45;
    wire logic g_2_45;
    assign p_2_45 = p_1_45 & p_1_43;
    assign g_2_45 = (p_1_45 & g_1_43) | g_1_45;
    wire logic p_2_47;
    wire logic g_2_47;
    assign p_2_47 = p_1_47 & p_1_45;
    assign g_2_47 = (p_1_47 & g_1_45) | g_1_47;
    wire logic p_2_49;
    wire logic g_2_49;
    assign p_2_49 = p_1_49 & p_1_47;
    assign g_2_49 = (p_1_49 & g_1_47) | g_1_49;
    wire logic p_2_51;
    wire logic g_2_51;
    assign p_2_51 = p_1_51 & p_1_49;
    assign g_2_51 = (p_1_51 & g_1_49) | g_1_51;
    wire logic p_2_53;
    wire logic g_2_53;
    assign p_2_53 = p_1_53 & p_1_51;
    assign g_2_53 = (p_1_53 & g_1_51) | g_1_53;
    wire logic p_2_55;
    wire logic g_2_55;
    assign p_2_55 = p_1_55 & p_1_53;
    assign g_2_55 = (p_1_55 & g_1_53) | g_1_55;
    wire logic p_2_57;
    wire logic g_2_57;
    assign p_2_57 = p_1_57 & p_1_55;
    assign g_2_57 = (p_1_57 & g_1_55) | g_1_57;
    wire logic p_2_59;
    wire logic g_2_59;
    assign p_2_59 = p_1_59 & p_1_57;
    assign g_2_59 = (p_1_59 & g_1_57) | g_1_59;
    wire logic p_2_61;
    wire logic g_2_61;
    assign p_2_61 = p_1_61 & p_1_59;
    assign g_2_61 = (p_1_61 & g_1_59) | g_1_61;
    wire logic p_2_63;
    wire logic g_2_63;
    assign p_2_63 = p_1_63 & p_1_61;
    assign g_2_63 = (p_1_63 & g_1_61) | g_1_63;
    wire logic p_2_65;
    wire logic g_2_65;
    assign p_2_65 = p_1_65 & p_1_63;
    assign g_2_65 = (p_1_65 & g_1_63) | g_1_65;
    wire logic p_2_67;
    wire logic g_2_67;
    assign p_2_67 = p_1_67 & p_1_65;
    assign g_2_67 = (p_1_67 & g_1_65) | g_1_67;
    wire logic p_2_69;
    wire logic g_2_69;
    assign p_2_69 = p_1_69 & p_1_67;
    assign g_2_69 = (p_1_69 & g_1_67) | g_1_69;
    wire logic p_2_71;
    wire logic g_2_71;
    assign p_2_71 = p_1_71 & p_1_69;
    assign g_2_71 = (p_1_71 & g_1_69) | g_1_71;
    wire logic p_2_73;
    wire logic g_2_73;
    assign p_2_73 = p_1_73 & p_1_71;
    assign g_2_73 = (p_1_73 & g_1_71) | g_1_73;
    wire logic p_2_75;
    wire logic g_2_75;
    assign p_2_75 = p_1_75 & p_1_73;
    assign g_2_75 = (p_1_75 & g_1_73) | g_1_75;
    wire logic p_2_77;
    wire logic g_2_77;
    assign p_2_77 = p_1_77 & p_1_75;
    assign g_2_77 = (p_1_77 & g_1_75) | g_1_77;
    wire logic p_2_79;
    wire logic g_2_79;
    assign p_2_79 = p_1_79 & p_1_77;
    assign g_2_79 = (p_1_79 & g_1_77) | g_1_79;
    wire logic p_2_81;
    wire logic g_2_81;
    assign p_2_81 = p_1_81 & p_1_79;
    assign g_2_81 = (p_1_81 & g_1_79) | g_1_81;
    wire logic p_2_83;
    wire logic g_2_83;
    assign p_2_83 = p_1_83 & p_1_81;
    assign g_2_83 = (p_1_83 & g_1_81) | g_1_83;
    wire logic p_2_85;
    wire logic g_2_85;
    assign p_2_85 = p_1_85 & p_1_83;
    assign g_2_85 = (p_1_85 & g_1_83) | g_1_85;
    wire logic p_2_87;
    wire logic g_2_87;
    assign p_2_87 = p_1_87 & p_1_85;
    assign g_2_87 = (p_1_87 & g_1_85) | g_1_87;
    wire logic p_2_89;
    wire logic g_2_89;
    assign p_2_89 = p_1_89 & p_1_87;
    assign g_2_89 = (p_1_89 & g_1_87) | g_1_89;
    wire logic p_2_91;
    wire logic g_2_91;
    assign p_2_91 = p_1_91 & p_1_89;
    assign g_2_91 = (p_1_91 & g_1_89) | g_1_91;
    wire logic p_2_93;
    wire logic g_2_93;
    assign p_2_93 = p_1_93 & p_1_91;
    assign g_2_93 = (p_1_93 & g_1_91) | g_1_93;
    wire logic p_2_95;
    wire logic g_2_95;
    assign p_2_95 = p_1_95 & p_1_93;
    assign g_2_95 = (p_1_95 & g_1_93) | g_1_95;
    wire logic p_2_97;
    wire logic g_2_97;
    assign p_2_97 = p_1_97 & p_1_95;
    assign g_2_97 = (p_1_97 & g_1_95) | g_1_97;
    wire logic p_2_99;
    wire logic g_2_99;
    assign p_2_99 = p_1_99 & p_1_97;
    assign g_2_99 = (p_1_99 & g_1_97) | g_1_99;
    wire logic p_2_101;
    wire logic g_2_101;
    assign p_2_101 = p_1_101 & p_1_99;
    assign g_2_101 = (p_1_101 & g_1_99) | g_1_101;
    wire logic p_2_103;
    wire logic g_2_103;
    assign p_2_103 = p_1_103 & p_1_101;
    assign g_2_103 = (p_1_103 & g_1_101) | g_1_103;
    wire logic p_2_105;
    wire logic g_2_105;
    assign p_2_105 = p_1_105 & p_1_103;
    assign g_2_105 = (p_1_105 & g_1_103) | g_1_105;
    wire logic p_2_107;
    wire logic g_2_107;
    assign p_2_107 = p_1_107 & p_1_105;
    assign g_2_107 = (p_1_107 & g_1_105) | g_1_107;
    wire logic p_2_109;
    wire logic g_2_109;
    assign p_2_109 = p_1_109 & p_1_107;
    assign g_2_109 = (p_1_109 & g_1_107) | g_1_109;
    wire logic p_2_111;
    wire logic g_2_111;
    assign p_2_111 = p_1_111 & p_1_109;
    assign g_2_111 = (p_1_111 & g_1_109) | g_1_111;
    wire logic p_2_113;
    wire logic g_2_113;
    assign p_2_113 = p_1_113 & p_1_111;
    assign g_2_113 = (p_1_113 & g_1_111) | g_1_113;
    wire logic p_2_115;
    wire logic g_2_115;
    assign p_2_115 = p_1_115 & p_1_113;
    assign g_2_115 = (p_1_115 & g_1_113) | g_1_115;
    wire logic p_2_117;
    wire logic g_2_117;
    assign p_2_117 = p_1_117 & p_1_115;
    assign g_2_117 = (p_1_117 & g_1_115) | g_1_117;
    wire logic p_2_119;
    wire logic g_2_119;
    assign p_2_119 = p_1_119 & p_1_117;
    assign g_2_119 = (p_1_119 & g_1_117) | g_1_119;
    wire logic p_2_121;
    wire logic g_2_121;
    assign p_2_121 = p_1_121 & p_1_119;
    assign g_2_121 = (p_1_121 & g_1_119) | g_1_121;
    wire logic p_2_123;
    wire logic g_2_123;
    assign p_2_123 = p_1_123 & p_1_121;
    assign g_2_123 = (p_1_123 & g_1_121) | g_1_123;
    wire logic p_2_125;
    wire logic g_2_125;
    assign p_2_125 = p_1_125 & p_1_123;
    assign g_2_125 = (p_1_125 & g_1_123) | g_1_125;
    wire logic p_2_127;
    wire logic g_2_127;
    assign p_2_127 = p_1_127 & p_1_125;
    assign g_2_127 = (p_1_127 & g_1_125) | g_1_127;
    
    // HC stage 3
    wire logic p_3_5;
    wire logic g_3_5;
    assign p_3_5 = p_2_5 & p_1_1;
    assign g_3_5 = (p_2_5 & g_1_1) | g_2_5;
    wire logic p_3_7;
    wire logic g_3_7;
    assign p_3_7 = p_2_7 & p_2_3;
    assign g_3_7 = (p_2_7 & g_2_3) | g_2_7;
    wire logic p_3_9;
    wire logic g_3_9;
    assign p_3_9 = p_2_9 & p_2_5;
    assign g_3_9 = (p_2_9 & g_2_5) | g_2_9;
    wire logic p_3_11;
    wire logic g_3_11;
    assign p_3_11 = p_2_11 & p_2_7;
    assign g_3_11 = (p_2_11 & g_2_7) | g_2_11;
    wire logic p_3_13;
    wire logic g_3_13;
    assign p_3_13 = p_2_13 & p_2_9;
    assign g_3_13 = (p_2_13 & g_2_9) | g_2_13;
    wire logic p_3_15;
    wire logic g_3_15;
    assign p_3_15 = p_2_15 & p_2_11;
    assign g_3_15 = (p_2_15 & g_2_11) | g_2_15;
    wire logic p_3_17;
    wire logic g_3_17;
    assign p_3_17 = p_2_17 & p_2_13;
    assign g_3_17 = (p_2_17 & g_2_13) | g_2_17;
    wire logic p_3_19;
    wire logic g_3_19;
    assign p_3_19 = p_2_19 & p_2_15;
    assign g_3_19 = (p_2_19 & g_2_15) | g_2_19;
    wire logic p_3_21;
    wire logic g_3_21;
    assign p_3_21 = p_2_21 & p_2_17;
    assign g_3_21 = (p_2_21 & g_2_17) | g_2_21;
    wire logic p_3_23;
    wire logic g_3_23;
    assign p_3_23 = p_2_23 & p_2_19;
    assign g_3_23 = (p_2_23 & g_2_19) | g_2_23;
    wire logic p_3_25;
    wire logic g_3_25;
    assign p_3_25 = p_2_25 & p_2_21;
    assign g_3_25 = (p_2_25 & g_2_21) | g_2_25;
    wire logic p_3_27;
    wire logic g_3_27;
    assign p_3_27 = p_2_27 & p_2_23;
    assign g_3_27 = (p_2_27 & g_2_23) | g_2_27;
    wire logic p_3_29;
    wire logic g_3_29;
    assign p_3_29 = p_2_29 & p_2_25;
    assign g_3_29 = (p_2_29 & g_2_25) | g_2_29;
    wire logic p_3_31;
    wire logic g_3_31;
    assign p_3_31 = p_2_31 & p_2_27;
    assign g_3_31 = (p_2_31 & g_2_27) | g_2_31;
    wire logic p_3_33;
    wire logic g_3_33;
    assign p_3_33 = p_2_33 & p_2_29;
    assign g_3_33 = (p_2_33 & g_2_29) | g_2_33;
    wire logic p_3_35;
    wire logic g_3_35;
    assign p_3_35 = p_2_35 & p_2_31;
    assign g_3_35 = (p_2_35 & g_2_31) | g_2_35;
    wire logic p_3_37;
    wire logic g_3_37;
    assign p_3_37 = p_2_37 & p_2_33;
    assign g_3_37 = (p_2_37 & g_2_33) | g_2_37;
    wire logic p_3_39;
    wire logic g_3_39;
    assign p_3_39 = p_2_39 & p_2_35;
    assign g_3_39 = (p_2_39 & g_2_35) | g_2_39;
    wire logic p_3_41;
    wire logic g_3_41;
    assign p_3_41 = p_2_41 & p_2_37;
    assign g_3_41 = (p_2_41 & g_2_37) | g_2_41;
    wire logic p_3_43;
    wire logic g_3_43;
    assign p_3_43 = p_2_43 & p_2_39;
    assign g_3_43 = (p_2_43 & g_2_39) | g_2_43;
    wire logic p_3_45;
    wire logic g_3_45;
    assign p_3_45 = p_2_45 & p_2_41;
    assign g_3_45 = (p_2_45 & g_2_41) | g_2_45;
    wire logic p_3_47;
    wire logic g_3_47;
    assign p_3_47 = p_2_47 & p_2_43;
    assign g_3_47 = (p_2_47 & g_2_43) | g_2_47;
    wire logic p_3_49;
    wire logic g_3_49;
    assign p_3_49 = p_2_49 & p_2_45;
    assign g_3_49 = (p_2_49 & g_2_45) | g_2_49;
    wire logic p_3_51;
    wire logic g_3_51;
    assign p_3_51 = p_2_51 & p_2_47;
    assign g_3_51 = (p_2_51 & g_2_47) | g_2_51;
    wire logic p_3_53;
    wire logic g_3_53;
    assign p_3_53 = p_2_53 & p_2_49;
    assign g_3_53 = (p_2_53 & g_2_49) | g_2_53;
    wire logic p_3_55;
    wire logic g_3_55;
    assign p_3_55 = p_2_55 & p_2_51;
    assign g_3_55 = (p_2_55 & g_2_51) | g_2_55;
    wire logic p_3_57;
    wire logic g_3_57;
    assign p_3_57 = p_2_57 & p_2_53;
    assign g_3_57 = (p_2_57 & g_2_53) | g_2_57;
    wire logic p_3_59;
    wire logic g_3_59;
    assign p_3_59 = p_2_59 & p_2_55;
    assign g_3_59 = (p_2_59 & g_2_55) | g_2_59;
    wire logic p_3_61;
    wire logic g_3_61;
    assign p_3_61 = p_2_61 & p_2_57;
    assign g_3_61 = (p_2_61 & g_2_57) | g_2_61;
    wire logic p_3_63;
    wire logic g_3_63;
    assign p_3_63 = p_2_63 & p_2_59;
    assign g_3_63 = (p_2_63 & g_2_59) | g_2_63;
    wire logic p_3_65;
    wire logic g_3_65;
    assign p_3_65 = p_2_65 & p_2_61;
    assign g_3_65 = (p_2_65 & g_2_61) | g_2_65;
    wire logic p_3_67;
    wire logic g_3_67;
    assign p_3_67 = p_2_67 & p_2_63;
    assign g_3_67 = (p_2_67 & g_2_63) | g_2_67;
    wire logic p_3_69;
    wire logic g_3_69;
    assign p_3_69 = p_2_69 & p_2_65;
    assign g_3_69 = (p_2_69 & g_2_65) | g_2_69;
    wire logic p_3_71;
    wire logic g_3_71;
    assign p_3_71 = p_2_71 & p_2_67;
    assign g_3_71 = (p_2_71 & g_2_67) | g_2_71;
    wire logic p_3_73;
    wire logic g_3_73;
    assign p_3_73 = p_2_73 & p_2_69;
    assign g_3_73 = (p_2_73 & g_2_69) | g_2_73;
    wire logic p_3_75;
    wire logic g_3_75;
    assign p_3_75 = p_2_75 & p_2_71;
    assign g_3_75 = (p_2_75 & g_2_71) | g_2_75;
    wire logic p_3_77;
    wire logic g_3_77;
    assign p_3_77 = p_2_77 & p_2_73;
    assign g_3_77 = (p_2_77 & g_2_73) | g_2_77;
    wire logic p_3_79;
    wire logic g_3_79;
    assign p_3_79 = p_2_79 & p_2_75;
    assign g_3_79 = (p_2_79 & g_2_75) | g_2_79;
    wire logic p_3_81;
    wire logic g_3_81;
    assign p_3_81 = p_2_81 & p_2_77;
    assign g_3_81 = (p_2_81 & g_2_77) | g_2_81;
    wire logic p_3_83;
    wire logic g_3_83;
    assign p_3_83 = p_2_83 & p_2_79;
    assign g_3_83 = (p_2_83 & g_2_79) | g_2_83;
    wire logic p_3_85;
    wire logic g_3_85;
    assign p_3_85 = p_2_85 & p_2_81;
    assign g_3_85 = (p_2_85 & g_2_81) | g_2_85;
    wire logic p_3_87;
    wire logic g_3_87;
    assign p_3_87 = p_2_87 & p_2_83;
    assign g_3_87 = (p_2_87 & g_2_83) | g_2_87;
    wire logic p_3_89;
    wire logic g_3_89;
    assign p_3_89 = p_2_89 & p_2_85;
    assign g_3_89 = (p_2_89 & g_2_85) | g_2_89;
    wire logic p_3_91;
    wire logic g_3_91;
    assign p_3_91 = p_2_91 & p_2_87;
    assign g_3_91 = (p_2_91 & g_2_87) | g_2_91;
    wire logic p_3_93;
    wire logic g_3_93;
    assign p_3_93 = p_2_93 & p_2_89;
    assign g_3_93 = (p_2_93 & g_2_89) | g_2_93;
    wire logic p_3_95;
    wire logic g_3_95;
    assign p_3_95 = p_2_95 & p_2_91;
    assign g_3_95 = (p_2_95 & g_2_91) | g_2_95;
    wire logic p_3_97;
    wire logic g_3_97;
    assign p_3_97 = p_2_97 & p_2_93;
    assign g_3_97 = (p_2_97 & g_2_93) | g_2_97;
    wire logic p_3_99;
    wire logic g_3_99;
    assign p_3_99 = p_2_99 & p_2_95;
    assign g_3_99 = (p_2_99 & g_2_95) | g_2_99;
    wire logic p_3_101;
    wire logic g_3_101;
    assign p_3_101 = p_2_101 & p_2_97;
    assign g_3_101 = (p_2_101 & g_2_97) | g_2_101;
    wire logic p_3_103;
    wire logic g_3_103;
    assign p_3_103 = p_2_103 & p_2_99;
    assign g_3_103 = (p_2_103 & g_2_99) | g_2_103;
    wire logic p_3_105;
    wire logic g_3_105;
    assign p_3_105 = p_2_105 & p_2_101;
    assign g_3_105 = (p_2_105 & g_2_101) | g_2_105;
    wire logic p_3_107;
    wire logic g_3_107;
    assign p_3_107 = p_2_107 & p_2_103;
    assign g_3_107 = (p_2_107 & g_2_103) | g_2_107;
    wire logic p_3_109;
    wire logic g_3_109;
    assign p_3_109 = p_2_109 & p_2_105;
    assign g_3_109 = (p_2_109 & g_2_105) | g_2_109;
    wire logic p_3_111;
    wire logic g_3_111;
    assign p_3_111 = p_2_111 & p_2_107;
    assign g_3_111 = (p_2_111 & g_2_107) | g_2_111;
    wire logic p_3_113;
    wire logic g_3_113;
    assign p_3_113 = p_2_113 & p_2_109;
    assign g_3_113 = (p_2_113 & g_2_109) | g_2_113;
    wire logic p_3_115;
    wire logic g_3_115;
    assign p_3_115 = p_2_115 & p_2_111;
    assign g_3_115 = (p_2_115 & g_2_111) | g_2_115;
    wire logic p_3_117;
    wire logic g_3_117;
    assign p_3_117 = p_2_117 & p_2_113;
    assign g_3_117 = (p_2_117 & g_2_113) | g_2_117;
    wire logic p_3_119;
    wire logic g_3_119;
    assign p_3_119 = p_2_119 & p_2_115;
    assign g_3_119 = (p_2_119 & g_2_115) | g_2_119;
    wire logic p_3_121;
    wire logic g_3_121;
    assign p_3_121 = p_2_121 & p_2_117;
    assign g_3_121 = (p_2_121 & g_2_117) | g_2_121;
    wire logic p_3_123;
    wire logic g_3_123;
    assign p_3_123 = p_2_123 & p_2_119;
    assign g_3_123 = (p_2_123 & g_2_119) | g_2_123;
    wire logic p_3_125;
    wire logic g_3_125;
    assign p_3_125 = p_2_125 & p_2_121;
    assign g_3_125 = (p_2_125 & g_2_121) | g_2_125;
    wire logic p_3_127;
    wire logic g_3_127;
    assign p_3_127 = p_2_127 & p_2_123;
    assign g_3_127 = (p_2_127 & g_2_123) | g_2_127;
    
    // HC stage 4
    wire logic p_4_9;
    wire logic g_4_9;
    assign p_4_9 = p_3_9 & p_1_1;
    assign g_4_9 = (p_3_9 & g_1_1) | g_3_9;
    wire logic p_4_11;
    wire logic g_4_11;
    assign p_4_11 = p_3_11 & p_2_3;
    assign g_4_11 = (p_3_11 & g_2_3) | g_3_11;
    wire logic p_4_13;
    wire logic g_4_13;
    assign p_4_13 = p_3_13 & p_3_5;
    assign g_4_13 = (p_3_13 & g_3_5) | g_3_13;
    wire logic p_4_15;
    wire logic g_4_15;
    assign p_4_15 = p_3_15 & p_3_7;
    assign g_4_15 = (p_3_15 & g_3_7) | g_3_15;
    wire logic p_4_17;
    wire logic g_4_17;
    assign p_4_17 = p_3_17 & p_3_9;
    assign g_4_17 = (p_3_17 & g_3_9) | g_3_17;
    wire logic p_4_19;
    wire logic g_4_19;
    assign p_4_19 = p_3_19 & p_3_11;
    assign g_4_19 = (p_3_19 & g_3_11) | g_3_19;
    wire logic p_4_21;
    wire logic g_4_21;
    assign p_4_21 = p_3_21 & p_3_13;
    assign g_4_21 = (p_3_21 & g_3_13) | g_3_21;
    wire logic p_4_23;
    wire logic g_4_23;
    assign p_4_23 = p_3_23 & p_3_15;
    assign g_4_23 = (p_3_23 & g_3_15) | g_3_23;
    wire logic p_4_25;
    wire logic g_4_25;
    assign p_4_25 = p_3_25 & p_3_17;
    assign g_4_25 = (p_3_25 & g_3_17) | g_3_25;
    wire logic p_4_27;
    wire logic g_4_27;
    assign p_4_27 = p_3_27 & p_3_19;
    assign g_4_27 = (p_3_27 & g_3_19) | g_3_27;
    wire logic p_4_29;
    wire logic g_4_29;
    assign p_4_29 = p_3_29 & p_3_21;
    assign g_4_29 = (p_3_29 & g_3_21) | g_3_29;
    wire logic p_4_31;
    wire logic g_4_31;
    assign p_4_31 = p_3_31 & p_3_23;
    assign g_4_31 = (p_3_31 & g_3_23) | g_3_31;
    wire logic p_4_33;
    wire logic g_4_33;
    assign p_4_33 = p_3_33 & p_3_25;
    assign g_4_33 = (p_3_33 & g_3_25) | g_3_33;
    wire logic p_4_35;
    wire logic g_4_35;
    assign p_4_35 = p_3_35 & p_3_27;
    assign g_4_35 = (p_3_35 & g_3_27) | g_3_35;
    wire logic p_4_37;
    wire logic g_4_37;
    assign p_4_37 = p_3_37 & p_3_29;
    assign g_4_37 = (p_3_37 & g_3_29) | g_3_37;
    wire logic p_4_39;
    wire logic g_4_39;
    assign p_4_39 = p_3_39 & p_3_31;
    assign g_4_39 = (p_3_39 & g_3_31) | g_3_39;
    wire logic p_4_41;
    wire logic g_4_41;
    assign p_4_41 = p_3_41 & p_3_33;
    assign g_4_41 = (p_3_41 & g_3_33) | g_3_41;
    wire logic p_4_43;
    wire logic g_4_43;
    assign p_4_43 = p_3_43 & p_3_35;
    assign g_4_43 = (p_3_43 & g_3_35) | g_3_43;
    wire logic p_4_45;
    wire logic g_4_45;
    assign p_4_45 = p_3_45 & p_3_37;
    assign g_4_45 = (p_3_45 & g_3_37) | g_3_45;
    wire logic p_4_47;
    wire logic g_4_47;
    assign p_4_47 = p_3_47 & p_3_39;
    assign g_4_47 = (p_3_47 & g_3_39) | g_3_47;
    wire logic p_4_49;
    wire logic g_4_49;
    assign p_4_49 = p_3_49 & p_3_41;
    assign g_4_49 = (p_3_49 & g_3_41) | g_3_49;
    wire logic p_4_51;
    wire logic g_4_51;
    assign p_4_51 = p_3_51 & p_3_43;
    assign g_4_51 = (p_3_51 & g_3_43) | g_3_51;
    wire logic p_4_53;
    wire logic g_4_53;
    assign p_4_53 = p_3_53 & p_3_45;
    assign g_4_53 = (p_3_53 & g_3_45) | g_3_53;
    wire logic p_4_55;
    wire logic g_4_55;
    assign p_4_55 = p_3_55 & p_3_47;
    assign g_4_55 = (p_3_55 & g_3_47) | g_3_55;
    wire logic p_4_57;
    wire logic g_4_57;
    assign p_4_57 = p_3_57 & p_3_49;
    assign g_4_57 = (p_3_57 & g_3_49) | g_3_57;
    wire logic p_4_59;
    wire logic g_4_59;
    assign p_4_59 = p_3_59 & p_3_51;
    assign g_4_59 = (p_3_59 & g_3_51) | g_3_59;
    wire logic p_4_61;
    wire logic g_4_61;
    assign p_4_61 = p_3_61 & p_3_53;
    assign g_4_61 = (p_3_61 & g_3_53) | g_3_61;
    wire logic p_4_63;
    wire logic g_4_63;
    assign p_4_63 = p_3_63 & p_3_55;
    assign g_4_63 = (p_3_63 & g_3_55) | g_3_63;
    wire logic p_4_65;
    wire logic g_4_65;
    assign p_4_65 = p_3_65 & p_3_57;
    assign g_4_65 = (p_3_65 & g_3_57) | g_3_65;
    wire logic p_4_67;
    wire logic g_4_67;
    assign p_4_67 = p_3_67 & p_3_59;
    assign g_4_67 = (p_3_67 & g_3_59) | g_3_67;
    wire logic p_4_69;
    wire logic g_4_69;
    assign p_4_69 = p_3_69 & p_3_61;
    assign g_4_69 = (p_3_69 & g_3_61) | g_3_69;
    wire logic p_4_71;
    wire logic g_4_71;
    assign p_4_71 = p_3_71 & p_3_63;
    assign g_4_71 = (p_3_71 & g_3_63) | g_3_71;
    wire logic p_4_73;
    wire logic g_4_73;
    assign p_4_73 = p_3_73 & p_3_65;
    assign g_4_73 = (p_3_73 & g_3_65) | g_3_73;
    wire logic p_4_75;
    wire logic g_4_75;
    assign p_4_75 = p_3_75 & p_3_67;
    assign g_4_75 = (p_3_75 & g_3_67) | g_3_75;
    wire logic p_4_77;
    wire logic g_4_77;
    assign p_4_77 = p_3_77 & p_3_69;
    assign g_4_77 = (p_3_77 & g_3_69) | g_3_77;
    wire logic p_4_79;
    wire logic g_4_79;
    assign p_4_79 = p_3_79 & p_3_71;
    assign g_4_79 = (p_3_79 & g_3_71) | g_3_79;
    wire logic p_4_81;
    wire logic g_4_81;
    assign p_4_81 = p_3_81 & p_3_73;
    assign g_4_81 = (p_3_81 & g_3_73) | g_3_81;
    wire logic p_4_83;
    wire logic g_4_83;
    assign p_4_83 = p_3_83 & p_3_75;
    assign g_4_83 = (p_3_83 & g_3_75) | g_3_83;
    wire logic p_4_85;
    wire logic g_4_85;
    assign p_4_85 = p_3_85 & p_3_77;
    assign g_4_85 = (p_3_85 & g_3_77) | g_3_85;
    wire logic p_4_87;
    wire logic g_4_87;
    assign p_4_87 = p_3_87 & p_3_79;
    assign g_4_87 = (p_3_87 & g_3_79) | g_3_87;
    wire logic p_4_89;
    wire logic g_4_89;
    assign p_4_89 = p_3_89 & p_3_81;
    assign g_4_89 = (p_3_89 & g_3_81) | g_3_89;
    wire logic p_4_91;
    wire logic g_4_91;
    assign p_4_91 = p_3_91 & p_3_83;
    assign g_4_91 = (p_3_91 & g_3_83) | g_3_91;
    wire logic p_4_93;
    wire logic g_4_93;
    assign p_4_93 = p_3_93 & p_3_85;
    assign g_4_93 = (p_3_93 & g_3_85) | g_3_93;
    wire logic p_4_95;
    wire logic g_4_95;
    assign p_4_95 = p_3_95 & p_3_87;
    assign g_4_95 = (p_3_95 & g_3_87) | g_3_95;
    wire logic p_4_97;
    wire logic g_4_97;
    assign p_4_97 = p_3_97 & p_3_89;
    assign g_4_97 = (p_3_97 & g_3_89) | g_3_97;
    wire logic p_4_99;
    wire logic g_4_99;
    assign p_4_99 = p_3_99 & p_3_91;
    assign g_4_99 = (p_3_99 & g_3_91) | g_3_99;
    wire logic p_4_101;
    wire logic g_4_101;
    assign p_4_101 = p_3_101 & p_3_93;
    assign g_4_101 = (p_3_101 & g_3_93) | g_3_101;
    wire logic p_4_103;
    wire logic g_4_103;
    assign p_4_103 = p_3_103 & p_3_95;
    assign g_4_103 = (p_3_103 & g_3_95) | g_3_103;
    wire logic p_4_105;
    wire logic g_4_105;
    assign p_4_105 = p_3_105 & p_3_97;
    assign g_4_105 = (p_3_105 & g_3_97) | g_3_105;
    wire logic p_4_107;
    wire logic g_4_107;
    assign p_4_107 = p_3_107 & p_3_99;
    assign g_4_107 = (p_3_107 & g_3_99) | g_3_107;
    wire logic p_4_109;
    wire logic g_4_109;
    assign p_4_109 = p_3_109 & p_3_101;
    assign g_4_109 = (p_3_109 & g_3_101) | g_3_109;
    wire logic p_4_111;
    wire logic g_4_111;
    assign p_4_111 = p_3_111 & p_3_103;
    assign g_4_111 = (p_3_111 & g_3_103) | g_3_111;
    wire logic p_4_113;
    wire logic g_4_113;
    assign p_4_113 = p_3_113 & p_3_105;
    assign g_4_113 = (p_3_113 & g_3_105) | g_3_113;
    wire logic p_4_115;
    wire logic g_4_115;
    assign p_4_115 = p_3_115 & p_3_107;
    assign g_4_115 = (p_3_115 & g_3_107) | g_3_115;
    wire logic p_4_117;
    wire logic g_4_117;
    assign p_4_117 = p_3_117 & p_3_109;
    assign g_4_117 = (p_3_117 & g_3_109) | g_3_117;
    wire logic p_4_119;
    wire logic g_4_119;
    assign p_4_119 = p_3_119 & p_3_111;
    assign g_4_119 = (p_3_119 & g_3_111) | g_3_119;
    wire logic p_4_121;
    wire logic g_4_121;
    assign p_4_121 = p_3_121 & p_3_113;
    assign g_4_121 = (p_3_121 & g_3_113) | g_3_121;
    wire logic p_4_123;
    wire logic g_4_123;
    assign p_4_123 = p_3_123 & p_3_115;
    assign g_4_123 = (p_3_123 & g_3_115) | g_3_123;
    wire logic p_4_125;
    wire logic g_4_125;
    assign p_4_125 = p_3_125 & p_3_117;
    assign g_4_125 = (p_3_125 & g_3_117) | g_3_125;
    wire logic p_4_127;
    wire logic g_4_127;
    assign p_4_127 = p_3_127 & p_3_119;
    assign g_4_127 = (p_3_127 & g_3_119) | g_3_127;
    
    // HC stage 5
    wire logic p_5_17;
    wire logic g_5_17;
    assign p_5_17 = p_4_17 & p_1_1;
    assign g_5_17 = (p_4_17 & g_1_1) | g_4_17;
    wire logic p_5_19;
    wire logic g_5_19;
    assign p_5_19 = p_4_19 & p_2_3;
    assign g_5_19 = (p_4_19 & g_2_3) | g_4_19;
    wire logic p_5_21;
    wire logic g_5_21;
    assign p_5_21 = p_4_21 & p_3_5;
    assign g_5_21 = (p_4_21 & g_3_5) | g_4_21;
    wire logic p_5_23;
    wire logic g_5_23;
    assign p_5_23 = p_4_23 & p_3_7;
    assign g_5_23 = (p_4_23 & g_3_7) | g_4_23;
    wire logic p_5_25;
    wire logic g_5_25;
    assign p_5_25 = p_4_25 & p_4_9;
    assign g_5_25 = (p_4_25 & g_4_9) | g_4_25;
    wire logic p_5_27;
    wire logic g_5_27;
    assign p_5_27 = p_4_27 & p_4_11;
    assign g_5_27 = (p_4_27 & g_4_11) | g_4_27;
    wire logic p_5_29;
    wire logic g_5_29;
    assign p_5_29 = p_4_29 & p_4_13;
    assign g_5_29 = (p_4_29 & g_4_13) | g_4_29;
    wire logic p_5_31;
    wire logic g_5_31;
    assign p_5_31 = p_4_31 & p_4_15;
    assign g_5_31 = (p_4_31 & g_4_15) | g_4_31;
    wire logic p_5_33;
    wire logic g_5_33;
    assign p_5_33 = p_4_33 & p_4_17;
    assign g_5_33 = (p_4_33 & g_4_17) | g_4_33;
    wire logic p_5_35;
    wire logic g_5_35;
    assign p_5_35 = p_4_35 & p_4_19;
    assign g_5_35 = (p_4_35 & g_4_19) | g_4_35;
    wire logic p_5_37;
    wire logic g_5_37;
    assign p_5_37 = p_4_37 & p_4_21;
    assign g_5_37 = (p_4_37 & g_4_21) | g_4_37;
    wire logic p_5_39;
    wire logic g_5_39;
    assign p_5_39 = p_4_39 & p_4_23;
    assign g_5_39 = (p_4_39 & g_4_23) | g_4_39;
    wire logic p_5_41;
    wire logic g_5_41;
    assign p_5_41 = p_4_41 & p_4_25;
    assign g_5_41 = (p_4_41 & g_4_25) | g_4_41;
    wire logic p_5_43;
    wire logic g_5_43;
    assign p_5_43 = p_4_43 & p_4_27;
    assign g_5_43 = (p_4_43 & g_4_27) | g_4_43;
    wire logic p_5_45;
    wire logic g_5_45;
    assign p_5_45 = p_4_45 & p_4_29;
    assign g_5_45 = (p_4_45 & g_4_29) | g_4_45;
    wire logic p_5_47;
    wire logic g_5_47;
    assign p_5_47 = p_4_47 & p_4_31;
    assign g_5_47 = (p_4_47 & g_4_31) | g_4_47;
    wire logic p_5_49;
    wire logic g_5_49;
    assign p_5_49 = p_4_49 & p_4_33;
    assign g_5_49 = (p_4_49 & g_4_33) | g_4_49;
    wire logic p_5_51;
    wire logic g_5_51;
    assign p_5_51 = p_4_51 & p_4_35;
    assign g_5_51 = (p_4_51 & g_4_35) | g_4_51;
    wire logic p_5_53;
    wire logic g_5_53;
    assign p_5_53 = p_4_53 & p_4_37;
    assign g_5_53 = (p_4_53 & g_4_37) | g_4_53;
    wire logic p_5_55;
    wire logic g_5_55;
    assign p_5_55 = p_4_55 & p_4_39;
    assign g_5_55 = (p_4_55 & g_4_39) | g_4_55;
    wire logic p_5_57;
    wire logic g_5_57;
    assign p_5_57 = p_4_57 & p_4_41;
    assign g_5_57 = (p_4_57 & g_4_41) | g_4_57;
    wire logic p_5_59;
    wire logic g_5_59;
    assign p_5_59 = p_4_59 & p_4_43;
    assign g_5_59 = (p_4_59 & g_4_43) | g_4_59;
    wire logic p_5_61;
    wire logic g_5_61;
    assign p_5_61 = p_4_61 & p_4_45;
    assign g_5_61 = (p_4_61 & g_4_45) | g_4_61;
    wire logic p_5_63;
    wire logic g_5_63;
    assign p_5_63 = p_4_63 & p_4_47;
    assign g_5_63 = (p_4_63 & g_4_47) | g_4_63;
    wire logic p_5_65;
    wire logic g_5_65;
    assign p_5_65 = p_4_65 & p_4_49;
    assign g_5_65 = (p_4_65 & g_4_49) | g_4_65;
    wire logic p_5_67;
    wire logic g_5_67;
    assign p_5_67 = p_4_67 & p_4_51;
    assign g_5_67 = (p_4_67 & g_4_51) | g_4_67;
    wire logic p_5_69;
    wire logic g_5_69;
    assign p_5_69 = p_4_69 & p_4_53;
    assign g_5_69 = (p_4_69 & g_4_53) | g_4_69;
    wire logic p_5_71;
    wire logic g_5_71;
    assign p_5_71 = p_4_71 & p_4_55;
    assign g_5_71 = (p_4_71 & g_4_55) | g_4_71;
    wire logic p_5_73;
    wire logic g_5_73;
    assign p_5_73 = p_4_73 & p_4_57;
    assign g_5_73 = (p_4_73 & g_4_57) | g_4_73;
    wire logic p_5_75;
    wire logic g_5_75;
    assign p_5_75 = p_4_75 & p_4_59;
    assign g_5_75 = (p_4_75 & g_4_59) | g_4_75;
    wire logic p_5_77;
    wire logic g_5_77;
    assign p_5_77 = p_4_77 & p_4_61;
    assign g_5_77 = (p_4_77 & g_4_61) | g_4_77;
    wire logic p_5_79;
    wire logic g_5_79;
    assign p_5_79 = p_4_79 & p_4_63;
    assign g_5_79 = (p_4_79 & g_4_63) | g_4_79;
    wire logic p_5_81;
    wire logic g_5_81;
    assign p_5_81 = p_4_81 & p_4_65;
    assign g_5_81 = (p_4_81 & g_4_65) | g_4_81;
    wire logic p_5_83;
    wire logic g_5_83;
    assign p_5_83 = p_4_83 & p_4_67;
    assign g_5_83 = (p_4_83 & g_4_67) | g_4_83;
    wire logic p_5_85;
    wire logic g_5_85;
    assign p_5_85 = p_4_85 & p_4_69;
    assign g_5_85 = (p_4_85 & g_4_69) | g_4_85;
    wire logic p_5_87;
    wire logic g_5_87;
    assign p_5_87 = p_4_87 & p_4_71;
    assign g_5_87 = (p_4_87 & g_4_71) | g_4_87;
    wire logic p_5_89;
    wire logic g_5_89;
    assign p_5_89 = p_4_89 & p_4_73;
    assign g_5_89 = (p_4_89 & g_4_73) | g_4_89;
    wire logic p_5_91;
    wire logic g_5_91;
    assign p_5_91 = p_4_91 & p_4_75;
    assign g_5_91 = (p_4_91 & g_4_75) | g_4_91;
    wire logic p_5_93;
    wire logic g_5_93;
    assign p_5_93 = p_4_93 & p_4_77;
    assign g_5_93 = (p_4_93 & g_4_77) | g_4_93;
    wire logic p_5_95;
    wire logic g_5_95;
    assign p_5_95 = p_4_95 & p_4_79;
    assign g_5_95 = (p_4_95 & g_4_79) | g_4_95;
    wire logic p_5_97;
    wire logic g_5_97;
    assign p_5_97 = p_4_97 & p_4_81;
    assign g_5_97 = (p_4_97 & g_4_81) | g_4_97;
    wire logic p_5_99;
    wire logic g_5_99;
    assign p_5_99 = p_4_99 & p_4_83;
    assign g_5_99 = (p_4_99 & g_4_83) | g_4_99;
    wire logic p_5_101;
    wire logic g_5_101;
    assign p_5_101 = p_4_101 & p_4_85;
    assign g_5_101 = (p_4_101 & g_4_85) | g_4_101;
    wire logic p_5_103;
    wire logic g_5_103;
    assign p_5_103 = p_4_103 & p_4_87;
    assign g_5_103 = (p_4_103 & g_4_87) | g_4_103;
    wire logic p_5_105;
    wire logic g_5_105;
    assign p_5_105 = p_4_105 & p_4_89;
    assign g_5_105 = (p_4_105 & g_4_89) | g_4_105;
    wire logic p_5_107;
    wire logic g_5_107;
    assign p_5_107 = p_4_107 & p_4_91;
    assign g_5_107 = (p_4_107 & g_4_91) | g_4_107;
    wire logic p_5_109;
    wire logic g_5_109;
    assign p_5_109 = p_4_109 & p_4_93;
    assign g_5_109 = (p_4_109 & g_4_93) | g_4_109;
    wire logic p_5_111;
    wire logic g_5_111;
    assign p_5_111 = p_4_111 & p_4_95;
    assign g_5_111 = (p_4_111 & g_4_95) | g_4_111;
    wire logic p_5_113;
    wire logic g_5_113;
    assign p_5_113 = p_4_113 & p_4_97;
    assign g_5_113 = (p_4_113 & g_4_97) | g_4_113;
    wire logic p_5_115;
    wire logic g_5_115;
    assign p_5_115 = p_4_115 & p_4_99;
    assign g_5_115 = (p_4_115 & g_4_99) | g_4_115;
    wire logic p_5_117;
    wire logic g_5_117;
    assign p_5_117 = p_4_117 & p_4_101;
    assign g_5_117 = (p_4_117 & g_4_101) | g_4_117;
    wire logic p_5_119;
    wire logic g_5_119;
    assign p_5_119 = p_4_119 & p_4_103;
    assign g_5_119 = (p_4_119 & g_4_103) | g_4_119;
    wire logic p_5_121;
    wire logic g_5_121;
    assign p_5_121 = p_4_121 & p_4_105;
    assign g_5_121 = (p_4_121 & g_4_105) | g_4_121;
    wire logic p_5_123;
    wire logic g_5_123;
    assign p_5_123 = p_4_123 & p_4_107;
    assign g_5_123 = (p_4_123 & g_4_107) | g_4_123;
    wire logic p_5_125;
    wire logic g_5_125;
    assign p_5_125 = p_4_125 & p_4_109;
    assign g_5_125 = (p_4_125 & g_4_109) | g_4_125;
    wire logic p_5_127;
    wire logic g_5_127;
    assign p_5_127 = p_4_127 & p_4_111;
    assign g_5_127 = (p_4_127 & g_4_111) | g_4_127;
    
    // HC stage 6
    wire logic p_6_33;
    wire logic g_6_33;
    assign p_6_33 = p_5_33 & p_1_1;
    assign g_6_33 = (p_5_33 & g_1_1) | g_5_33;
    wire logic p_6_35;
    wire logic g_6_35;
    assign p_6_35 = p_5_35 & p_2_3;
    assign g_6_35 = (p_5_35 & g_2_3) | g_5_35;
    wire logic p_6_37;
    wire logic g_6_37;
    assign p_6_37 = p_5_37 & p_3_5;
    assign g_6_37 = (p_5_37 & g_3_5) | g_5_37;
    wire logic p_6_39;
    wire logic g_6_39;
    assign p_6_39 = p_5_39 & p_3_7;
    assign g_6_39 = (p_5_39 & g_3_7) | g_5_39;
    wire logic p_6_41;
    wire logic g_6_41;
    assign p_6_41 = p_5_41 & p_4_9;
    assign g_6_41 = (p_5_41 & g_4_9) | g_5_41;
    wire logic p_6_43;
    wire logic g_6_43;
    assign p_6_43 = p_5_43 & p_4_11;
    assign g_6_43 = (p_5_43 & g_4_11) | g_5_43;
    wire logic p_6_45;
    wire logic g_6_45;
    assign p_6_45 = p_5_45 & p_4_13;
    assign g_6_45 = (p_5_45 & g_4_13) | g_5_45;
    wire logic p_6_47;
    wire logic g_6_47;
    assign p_6_47 = p_5_47 & p_4_15;
    assign g_6_47 = (p_5_47 & g_4_15) | g_5_47;
    wire logic p_6_49;
    wire logic g_6_49;
    assign p_6_49 = p_5_49 & p_5_17;
    assign g_6_49 = (p_5_49 & g_5_17) | g_5_49;
    wire logic p_6_51;
    wire logic g_6_51;
    assign p_6_51 = p_5_51 & p_5_19;
    assign g_6_51 = (p_5_51 & g_5_19) | g_5_51;
    wire logic p_6_53;
    wire logic g_6_53;
    assign p_6_53 = p_5_53 & p_5_21;
    assign g_6_53 = (p_5_53 & g_5_21) | g_5_53;
    wire logic p_6_55;
    wire logic g_6_55;
    assign p_6_55 = p_5_55 & p_5_23;
    assign g_6_55 = (p_5_55 & g_5_23) | g_5_55;
    wire logic p_6_57;
    wire logic g_6_57;
    assign p_6_57 = p_5_57 & p_5_25;
    assign g_6_57 = (p_5_57 & g_5_25) | g_5_57;
    wire logic p_6_59;
    wire logic g_6_59;
    assign p_6_59 = p_5_59 & p_5_27;
    assign g_6_59 = (p_5_59 & g_5_27) | g_5_59;
    wire logic p_6_61;
    wire logic g_6_61;
    assign p_6_61 = p_5_61 & p_5_29;
    assign g_6_61 = (p_5_61 & g_5_29) | g_5_61;
    wire logic p_6_63;
    wire logic g_6_63;
    assign p_6_63 = p_5_63 & p_5_31;
    assign g_6_63 = (p_5_63 & g_5_31) | g_5_63;
    wire logic p_6_65;
    wire logic g_6_65;
    assign p_6_65 = p_5_65 & p_5_33;
    assign g_6_65 = (p_5_65 & g_5_33) | g_5_65;
    wire logic p_6_67;
    wire logic g_6_67;
    assign p_6_67 = p_5_67 & p_5_35;
    assign g_6_67 = (p_5_67 & g_5_35) | g_5_67;
    wire logic p_6_69;
    wire logic g_6_69;
    assign p_6_69 = p_5_69 & p_5_37;
    assign g_6_69 = (p_5_69 & g_5_37) | g_5_69;
    wire logic p_6_71;
    wire logic g_6_71;
    assign p_6_71 = p_5_71 & p_5_39;
    assign g_6_71 = (p_5_71 & g_5_39) | g_5_71;
    wire logic p_6_73;
    wire logic g_6_73;
    assign p_6_73 = p_5_73 & p_5_41;
    assign g_6_73 = (p_5_73 & g_5_41) | g_5_73;
    wire logic p_6_75;
    wire logic g_6_75;
    assign p_6_75 = p_5_75 & p_5_43;
    assign g_6_75 = (p_5_75 & g_5_43) | g_5_75;
    wire logic p_6_77;
    wire logic g_6_77;
    assign p_6_77 = p_5_77 & p_5_45;
    assign g_6_77 = (p_5_77 & g_5_45) | g_5_77;
    wire logic p_6_79;
    wire logic g_6_79;
    assign p_6_79 = p_5_79 & p_5_47;
    assign g_6_79 = (p_5_79 & g_5_47) | g_5_79;
    wire logic p_6_81;
    wire logic g_6_81;
    assign p_6_81 = p_5_81 & p_5_49;
    assign g_6_81 = (p_5_81 & g_5_49) | g_5_81;
    wire logic p_6_83;
    wire logic g_6_83;
    assign p_6_83 = p_5_83 & p_5_51;
    assign g_6_83 = (p_5_83 & g_5_51) | g_5_83;
    wire logic p_6_85;
    wire logic g_6_85;
    assign p_6_85 = p_5_85 & p_5_53;
    assign g_6_85 = (p_5_85 & g_5_53) | g_5_85;
    wire logic p_6_87;
    wire logic g_6_87;
    assign p_6_87 = p_5_87 & p_5_55;
    assign g_6_87 = (p_5_87 & g_5_55) | g_5_87;
    wire logic p_6_89;
    wire logic g_6_89;
    assign p_6_89 = p_5_89 & p_5_57;
    assign g_6_89 = (p_5_89 & g_5_57) | g_5_89;
    wire logic p_6_91;
    wire logic g_6_91;
    assign p_6_91 = p_5_91 & p_5_59;
    assign g_6_91 = (p_5_91 & g_5_59) | g_5_91;
    wire logic p_6_93;
    wire logic g_6_93;
    assign p_6_93 = p_5_93 & p_5_61;
    assign g_6_93 = (p_5_93 & g_5_61) | g_5_93;
    wire logic p_6_95;
    wire logic g_6_95;
    assign p_6_95 = p_5_95 & p_5_63;
    assign g_6_95 = (p_5_95 & g_5_63) | g_5_95;
    wire logic p_6_97;
    wire logic g_6_97;
    assign p_6_97 = p_5_97 & p_5_65;
    assign g_6_97 = (p_5_97 & g_5_65) | g_5_97;
    wire logic p_6_99;
    wire logic g_6_99;
    assign p_6_99 = p_5_99 & p_5_67;
    assign g_6_99 = (p_5_99 & g_5_67) | g_5_99;
    wire logic p_6_101;
    wire logic g_6_101;
    assign p_6_101 = p_5_101 & p_5_69;
    assign g_6_101 = (p_5_101 & g_5_69) | g_5_101;
    wire logic p_6_103;
    wire logic g_6_103;
    assign p_6_103 = p_5_103 & p_5_71;
    assign g_6_103 = (p_5_103 & g_5_71) | g_5_103;
    wire logic p_6_105;
    wire logic g_6_105;
    assign p_6_105 = p_5_105 & p_5_73;
    assign g_6_105 = (p_5_105 & g_5_73) | g_5_105;
    wire logic p_6_107;
    wire logic g_6_107;
    assign p_6_107 = p_5_107 & p_5_75;
    assign g_6_107 = (p_5_107 & g_5_75) | g_5_107;
    wire logic p_6_109;
    wire logic g_6_109;
    assign p_6_109 = p_5_109 & p_5_77;
    assign g_6_109 = (p_5_109 & g_5_77) | g_5_109;
    wire logic p_6_111;
    wire logic g_6_111;
    assign p_6_111 = p_5_111 & p_5_79;
    assign g_6_111 = (p_5_111 & g_5_79) | g_5_111;
    wire logic p_6_113;
    wire logic g_6_113;
    assign p_6_113 = p_5_113 & p_5_81;
    assign g_6_113 = (p_5_113 & g_5_81) | g_5_113;
    wire logic p_6_115;
    wire logic g_6_115;
    assign p_6_115 = p_5_115 & p_5_83;
    assign g_6_115 = (p_5_115 & g_5_83) | g_5_115;
    wire logic p_6_117;
    wire logic g_6_117;
    assign p_6_117 = p_5_117 & p_5_85;
    assign g_6_117 = (p_5_117 & g_5_85) | g_5_117;
    wire logic p_6_119;
    wire logic g_6_119;
    assign p_6_119 = p_5_119 & p_5_87;
    assign g_6_119 = (p_5_119 & g_5_87) | g_5_119;
    wire logic p_6_121;
    wire logic g_6_121;
    assign p_6_121 = p_5_121 & p_5_89;
    assign g_6_121 = (p_5_121 & g_5_89) | g_5_121;
    wire logic p_6_123;
    wire logic g_6_123;
    assign p_6_123 = p_5_123 & p_5_91;
    assign g_6_123 = (p_5_123 & g_5_91) | g_5_123;
    wire logic p_6_125;
    wire logic g_6_125;
    assign p_6_125 = p_5_125 & p_5_93;
    assign g_6_125 = (p_5_125 & g_5_93) | g_5_125;
    wire logic p_6_127;
    wire logic g_6_127;
    assign p_6_127 = p_5_127 & p_5_95;
    assign g_6_127 = (p_5_127 & g_5_95) | g_5_127;
    
    // HC stage 7
    wire logic p_7_65;
    wire logic g_7_65;
    assign p_7_65 = p_6_65 & p_1_1;
    assign g_7_65 = (p_6_65 & g_1_1) | g_6_65;
    wire logic p_7_67;
    wire logic g_7_67;
    assign p_7_67 = p_6_67 & p_2_3;
    assign g_7_67 = (p_6_67 & g_2_3) | g_6_67;
    wire logic p_7_69;
    wire logic g_7_69;
    assign p_7_69 = p_6_69 & p_3_5;
    assign g_7_69 = (p_6_69 & g_3_5) | g_6_69;
    wire logic p_7_71;
    wire logic g_7_71;
    assign p_7_71 = p_6_71 & p_3_7;
    assign g_7_71 = (p_6_71 & g_3_7) | g_6_71;
    wire logic p_7_73;
    wire logic g_7_73;
    assign p_7_73 = p_6_73 & p_4_9;
    assign g_7_73 = (p_6_73 & g_4_9) | g_6_73;
    wire logic p_7_75;
    wire logic g_7_75;
    assign p_7_75 = p_6_75 & p_4_11;
    assign g_7_75 = (p_6_75 & g_4_11) | g_6_75;
    wire logic p_7_77;
    wire logic g_7_77;
    assign p_7_77 = p_6_77 & p_4_13;
    assign g_7_77 = (p_6_77 & g_4_13) | g_6_77;
    wire logic p_7_79;
    wire logic g_7_79;
    assign p_7_79 = p_6_79 & p_4_15;
    assign g_7_79 = (p_6_79 & g_4_15) | g_6_79;
    wire logic p_7_81;
    wire logic g_7_81;
    assign p_7_81 = p_6_81 & p_5_17;
    assign g_7_81 = (p_6_81 & g_5_17) | g_6_81;
    wire logic p_7_83;
    wire logic g_7_83;
    assign p_7_83 = p_6_83 & p_5_19;
    assign g_7_83 = (p_6_83 & g_5_19) | g_6_83;
    wire logic p_7_85;
    wire logic g_7_85;
    assign p_7_85 = p_6_85 & p_5_21;
    assign g_7_85 = (p_6_85 & g_5_21) | g_6_85;
    wire logic p_7_87;
    wire logic g_7_87;
    assign p_7_87 = p_6_87 & p_5_23;
    assign g_7_87 = (p_6_87 & g_5_23) | g_6_87;
    wire logic p_7_89;
    wire logic g_7_89;
    assign p_7_89 = p_6_89 & p_5_25;
    assign g_7_89 = (p_6_89 & g_5_25) | g_6_89;
    wire logic p_7_91;
    wire logic g_7_91;
    assign p_7_91 = p_6_91 & p_5_27;
    assign g_7_91 = (p_6_91 & g_5_27) | g_6_91;
    wire logic p_7_93;
    wire logic g_7_93;
    assign p_7_93 = p_6_93 & p_5_29;
    assign g_7_93 = (p_6_93 & g_5_29) | g_6_93;
    wire logic p_7_95;
    wire logic g_7_95;
    assign p_7_95 = p_6_95 & p_5_31;
    assign g_7_95 = (p_6_95 & g_5_31) | g_6_95;
    wire logic p_7_97;
    wire logic g_7_97;
    assign p_7_97 = p_6_97 & p_6_33;
    assign g_7_97 = (p_6_97 & g_6_33) | g_6_97;
    wire logic p_7_99;
    wire logic g_7_99;
    assign p_7_99 = p_6_99 & p_6_35;
    assign g_7_99 = (p_6_99 & g_6_35) | g_6_99;
    wire logic p_7_101;
    wire logic g_7_101;
    assign p_7_101 = p_6_101 & p_6_37;
    assign g_7_101 = (p_6_101 & g_6_37) | g_6_101;
    wire logic p_7_103;
    wire logic g_7_103;
    assign p_7_103 = p_6_103 & p_6_39;
    assign g_7_103 = (p_6_103 & g_6_39) | g_6_103;
    wire logic p_7_105;
    wire logic g_7_105;
    assign p_7_105 = p_6_105 & p_6_41;
    assign g_7_105 = (p_6_105 & g_6_41) | g_6_105;
    wire logic p_7_107;
    wire logic g_7_107;
    assign p_7_107 = p_6_107 & p_6_43;
    assign g_7_107 = (p_6_107 & g_6_43) | g_6_107;
    wire logic p_7_109;
    wire logic g_7_109;
    assign p_7_109 = p_6_109 & p_6_45;
    assign g_7_109 = (p_6_109 & g_6_45) | g_6_109;
    wire logic p_7_111;
    wire logic g_7_111;
    assign p_7_111 = p_6_111 & p_6_47;
    assign g_7_111 = (p_6_111 & g_6_47) | g_6_111;
    wire logic p_7_113;
    wire logic g_7_113;
    assign p_7_113 = p_6_113 & p_6_49;
    assign g_7_113 = (p_6_113 & g_6_49) | g_6_113;
    wire logic p_7_115;
    wire logic g_7_115;
    assign p_7_115 = p_6_115 & p_6_51;
    assign g_7_115 = (p_6_115 & g_6_51) | g_6_115;
    wire logic p_7_117;
    wire logic g_7_117;
    assign p_7_117 = p_6_117 & p_6_53;
    assign g_7_117 = (p_6_117 & g_6_53) | g_6_117;
    wire logic p_7_119;
    wire logic g_7_119;
    assign p_7_119 = p_6_119 & p_6_55;
    assign g_7_119 = (p_6_119 & g_6_55) | g_6_119;
    wire logic p_7_121;
    wire logic g_7_121;
    assign p_7_121 = p_6_121 & p_6_57;
    assign g_7_121 = (p_6_121 & g_6_57) | g_6_121;
    wire logic p_7_123;
    wire logic g_7_123;
    assign p_7_123 = p_6_123 & p_6_59;
    assign g_7_123 = (p_6_123 & g_6_59) | g_6_123;
    wire logic p_7_125;
    wire logic g_7_125;
    assign p_7_125 = p_6_125 & p_6_61;
    assign g_7_125 = (p_6_125 & g_6_61) | g_6_125;
    wire logic p_7_127;
    wire logic g_7_127;
    assign p_7_127 = p_6_127 & p_6_63;
    assign g_7_127 = (p_6_127 & g_6_63) | g_6_127;
    
    // HC stage 8
    wire logic p_8_2;
    wire logic g_8_2;
    assign p_8_2 = p_0[2] & p_1_1;
    assign g_8_2 = (p_0[2] & g_1_1) | g_0[2];
    wire logic p_8_4;
    wire logic g_8_4;
    assign p_8_4 = p_0[4] & p_2_3;
    assign g_8_4 = (p_0[4] & g_2_3) | g_0[4];
    wire logic p_8_6;
    wire logic g_8_6;
    assign p_8_6 = p_0[6] & p_3_5;
    assign g_8_6 = (p_0[6] & g_3_5) | g_0[6];
    wire logic p_8_8;
    wire logic g_8_8;
    assign p_8_8 = p_0[8] & p_3_7;
    assign g_8_8 = (p_0[8] & g_3_7) | g_0[8];
    wire logic p_8_10;
    wire logic g_8_10;
    assign p_8_10 = p_0[10] & p_4_9;
    assign g_8_10 = (p_0[10] & g_4_9) | g_0[10];
    wire logic p_8_12;
    wire logic g_8_12;
    assign p_8_12 = p_0[12] & p_4_11;
    assign g_8_12 = (p_0[12] & g_4_11) | g_0[12];
    wire logic p_8_14;
    wire logic g_8_14;
    assign p_8_14 = p_0[14] & p_4_13;
    assign g_8_14 = (p_0[14] & g_4_13) | g_0[14];
    wire logic p_8_16;
    wire logic g_8_16;
    assign p_8_16 = p_0[16] & p_4_15;
    assign g_8_16 = (p_0[16] & g_4_15) | g_0[16];
    wire logic p_8_18;
    wire logic g_8_18;
    assign p_8_18 = p_0[18] & p_5_17;
    assign g_8_18 = (p_0[18] & g_5_17) | g_0[18];
    wire logic p_8_20;
    wire logic g_8_20;
    assign p_8_20 = p_0[20] & p_5_19;
    assign g_8_20 = (p_0[20] & g_5_19) | g_0[20];
    wire logic p_8_22;
    wire logic g_8_22;
    assign p_8_22 = p_0[22] & p_5_21;
    assign g_8_22 = (p_0[22] & g_5_21) | g_0[22];
    wire logic p_8_24;
    wire logic g_8_24;
    assign p_8_24 = p_0[24] & p_5_23;
    assign g_8_24 = (p_0[24] & g_5_23) | g_0[24];
    wire logic p_8_26;
    wire logic g_8_26;
    assign p_8_26 = p_0[26] & p_5_25;
    assign g_8_26 = (p_0[26] & g_5_25) | g_0[26];
    wire logic p_8_28;
    wire logic g_8_28;
    assign p_8_28 = p_0[28] & p_5_27;
    assign g_8_28 = (p_0[28] & g_5_27) | g_0[28];
    wire logic p_8_30;
    wire logic g_8_30;
    assign p_8_30 = p_0[30] & p_5_29;
    assign g_8_30 = (p_0[30] & g_5_29) | g_0[30];
    wire logic p_8_32;
    wire logic g_8_32;
    assign p_8_32 = p_0[32] & p_5_31;
    assign g_8_32 = (p_0[32] & g_5_31) | g_0[32];
    wire logic p_8_34;
    wire logic g_8_34;
    assign p_8_34 = p_0[34] & p_6_33;
    assign g_8_34 = (p_0[34] & g_6_33) | g_0[34];
    wire logic p_8_36;
    wire logic g_8_36;
    assign p_8_36 = p_0[36] & p_6_35;
    assign g_8_36 = (p_0[36] & g_6_35) | g_0[36];
    wire logic p_8_38;
    wire logic g_8_38;
    assign p_8_38 = p_0[38] & p_6_37;
    assign g_8_38 = (p_0[38] & g_6_37) | g_0[38];
    wire logic p_8_40;
    wire logic g_8_40;
    assign p_8_40 = p_0[40] & p_6_39;
    assign g_8_40 = (p_0[40] & g_6_39) | g_0[40];
    wire logic p_8_42;
    wire logic g_8_42;
    assign p_8_42 = p_0[42] & p_6_41;
    assign g_8_42 = (p_0[42] & g_6_41) | g_0[42];
    wire logic p_8_44;
    wire logic g_8_44;
    assign p_8_44 = p_0[44] & p_6_43;
    assign g_8_44 = (p_0[44] & g_6_43) | g_0[44];
    wire logic p_8_46;
    wire logic g_8_46;
    assign p_8_46 = p_0[46] & p_6_45;
    assign g_8_46 = (p_0[46] & g_6_45) | g_0[46];
    wire logic p_8_48;
    wire logic g_8_48;
    assign p_8_48 = p_0[48] & p_6_47;
    assign g_8_48 = (p_0[48] & g_6_47) | g_0[48];
    wire logic p_8_50;
    wire logic g_8_50;
    assign p_8_50 = p_0[50] & p_6_49;
    assign g_8_50 = (p_0[50] & g_6_49) | g_0[50];
    wire logic p_8_52;
    wire logic g_8_52;
    assign p_8_52 = p_0[52] & p_6_51;
    assign g_8_52 = (p_0[52] & g_6_51) | g_0[52];
    wire logic p_8_54;
    wire logic g_8_54;
    assign p_8_54 = p_0[54] & p_6_53;
    assign g_8_54 = (p_0[54] & g_6_53) | g_0[54];
    wire logic p_8_56;
    wire logic g_8_56;
    assign p_8_56 = p_0[56] & p_6_55;
    assign g_8_56 = (p_0[56] & g_6_55) | g_0[56];
    wire logic p_8_58;
    wire logic g_8_58;
    assign p_8_58 = p_0[58] & p_6_57;
    assign g_8_58 = (p_0[58] & g_6_57) | g_0[58];
    wire logic p_8_60;
    wire logic g_8_60;
    assign p_8_60 = p_0[60] & p_6_59;
    assign g_8_60 = (p_0[60] & g_6_59) | g_0[60];
    wire logic p_8_62;
    wire logic g_8_62;
    assign p_8_62 = p_0[62] & p_6_61;
    assign g_8_62 = (p_0[62] & g_6_61) | g_0[62];
    wire logic p_8_64;
    wire logic g_8_64;
    assign p_8_64 = p_0[64] & p_6_63;
    assign g_8_64 = (p_0[64] & g_6_63) | g_0[64];
    wire logic p_8_66;
    wire logic g_8_66;
    assign p_8_66 = p_0[66] & p_7_65;
    assign g_8_66 = (p_0[66] & g_7_65) | g_0[66];
    wire logic p_8_68;
    wire logic g_8_68;
    assign p_8_68 = p_0[68] & p_7_67;
    assign g_8_68 = (p_0[68] & g_7_67) | g_0[68];
    wire logic p_8_70;
    wire logic g_8_70;
    assign p_8_70 = p_0[70] & p_7_69;
    assign g_8_70 = (p_0[70] & g_7_69) | g_0[70];
    wire logic p_8_72;
    wire logic g_8_72;
    assign p_8_72 = p_0[72] & p_7_71;
    assign g_8_72 = (p_0[72] & g_7_71) | g_0[72];
    wire logic p_8_74;
    wire logic g_8_74;
    assign p_8_74 = p_0[74] & p_7_73;
    assign g_8_74 = (p_0[74] & g_7_73) | g_0[74];
    wire logic p_8_76;
    wire logic g_8_76;
    assign p_8_76 = p_0[76] & p_7_75;
    assign g_8_76 = (p_0[76] & g_7_75) | g_0[76];
    wire logic p_8_78;
    wire logic g_8_78;
    assign p_8_78 = p_0[78] & p_7_77;
    assign g_8_78 = (p_0[78] & g_7_77) | g_0[78];
    wire logic p_8_80;
    wire logic g_8_80;
    assign p_8_80 = p_0[80] & p_7_79;
    assign g_8_80 = (p_0[80] & g_7_79) | g_0[80];
    wire logic p_8_82;
    wire logic g_8_82;
    assign p_8_82 = p_0[82] & p_7_81;
    assign g_8_82 = (p_0[82] & g_7_81) | g_0[82];
    wire logic p_8_84;
    wire logic g_8_84;
    assign p_8_84 = p_0[84] & p_7_83;
    assign g_8_84 = (p_0[84] & g_7_83) | g_0[84];
    wire logic p_8_86;
    wire logic g_8_86;
    assign p_8_86 = p_0[86] & p_7_85;
    assign g_8_86 = (p_0[86] & g_7_85) | g_0[86];
    wire logic p_8_88;
    wire logic g_8_88;
    assign p_8_88 = p_0[88] & p_7_87;
    assign g_8_88 = (p_0[88] & g_7_87) | g_0[88];
    wire logic p_8_90;
    wire logic g_8_90;
    assign p_8_90 = p_0[90] & p_7_89;
    assign g_8_90 = (p_0[90] & g_7_89) | g_0[90];
    wire logic p_8_92;
    wire logic g_8_92;
    assign p_8_92 = p_0[92] & p_7_91;
    assign g_8_92 = (p_0[92] & g_7_91) | g_0[92];
    wire logic p_8_94;
    wire logic g_8_94;
    assign p_8_94 = p_0[94] & p_7_93;
    assign g_8_94 = (p_0[94] & g_7_93) | g_0[94];
    wire logic p_8_96;
    wire logic g_8_96;
    assign p_8_96 = p_0[96] & p_7_95;
    assign g_8_96 = (p_0[96] & g_7_95) | g_0[96];
    wire logic p_8_98;
    wire logic g_8_98;
    assign p_8_98 = p_0[98] & p_7_97;
    assign g_8_98 = (p_0[98] & g_7_97) | g_0[98];
    wire logic p_8_100;
    wire logic g_8_100;
    assign p_8_100 = p_0[100] & p_7_99;
    assign g_8_100 = (p_0[100] & g_7_99) | g_0[100];
    wire logic p_8_102;
    wire logic g_8_102;
    assign p_8_102 = p_0[102] & p_7_101;
    assign g_8_102 = (p_0[102] & g_7_101) | g_0[102];
    wire logic p_8_104;
    wire logic g_8_104;
    assign p_8_104 = p_0[104] & p_7_103;
    assign g_8_104 = (p_0[104] & g_7_103) | g_0[104];
    wire logic p_8_106;
    wire logic g_8_106;
    assign p_8_106 = p_0[106] & p_7_105;
    assign g_8_106 = (p_0[106] & g_7_105) | g_0[106];
    wire logic p_8_108;
    wire logic g_8_108;
    assign p_8_108 = p_0[108] & p_7_107;
    assign g_8_108 = (p_0[108] & g_7_107) | g_0[108];
    wire logic p_8_110;
    wire logic g_8_110;
    assign p_8_110 = p_0[110] & p_7_109;
    assign g_8_110 = (p_0[110] & g_7_109) | g_0[110];
    wire logic p_8_112;
    wire logic g_8_112;
    assign p_8_112 = p_0[112] & p_7_111;
    assign g_8_112 = (p_0[112] & g_7_111) | g_0[112];
    wire logic p_8_114;
    wire logic g_8_114;
    assign p_8_114 = p_0[114] & p_7_113;
    assign g_8_114 = (p_0[114] & g_7_113) | g_0[114];
    wire logic p_8_116;
    wire logic g_8_116;
    assign p_8_116 = p_0[116] & p_7_115;
    assign g_8_116 = (p_0[116] & g_7_115) | g_0[116];
    wire logic p_8_118;
    wire logic g_8_118;
    assign p_8_118 = p_0[118] & p_7_117;
    assign g_8_118 = (p_0[118] & g_7_117) | g_0[118];
    wire logic p_8_120;
    wire logic g_8_120;
    assign p_8_120 = p_0[120] & p_7_119;
    assign g_8_120 = (p_0[120] & g_7_119) | g_0[120];
    wire logic p_8_122;
    wire logic g_8_122;
    assign p_8_122 = p_0[122] & p_7_121;
    assign g_8_122 = (p_0[122] & g_7_121) | g_0[122];
    wire logic p_8_124;
    wire logic g_8_124;
    assign p_8_124 = p_0[124] & p_7_123;
    assign g_8_124 = (p_0[124] & g_7_123) | g_0[124];
    wire logic p_8_126;
    wire logic g_8_126;
    assign p_8_126 = p_0[126] & p_7_125;
    assign g_8_126 = (p_0[126] & g_7_125) | g_0[126];
    
    // HC postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = p_0[3] ^ g_8_2;
    assign OUT[4] = p_0[4] ^ g_2_3;
    assign OUT[5] = p_0[5] ^ g_8_4;
    assign OUT[6] = p_0[6] ^ g_3_5;
    assign OUT[7] = p_0[7] ^ g_8_6;
    assign OUT[8] = p_0[8] ^ g_3_7;
    assign OUT[9] = p_0[9] ^ g_8_8;
    assign OUT[10] = p_0[10] ^ g_4_9;
    assign OUT[11] = p_0[11] ^ g_8_10;
    assign OUT[12] = p_0[12] ^ g_4_11;
    assign OUT[13] = p_0[13] ^ g_8_12;
    assign OUT[14] = p_0[14] ^ g_4_13;
    assign OUT[15] = p_0[15] ^ g_8_14;
    assign OUT[16] = p_0[16] ^ g_4_15;
    assign OUT[17] = p_0[17] ^ g_8_16;
    assign OUT[18] = p_0[18] ^ g_5_17;
    assign OUT[19] = p_0[19] ^ g_8_18;
    assign OUT[20] = p_0[20] ^ g_5_19;
    assign OUT[21] = p_0[21] ^ g_8_20;
    assign OUT[22] = p_0[22] ^ g_5_21;
    assign OUT[23] = p_0[23] ^ g_8_22;
    assign OUT[24] = p_0[24] ^ g_5_23;
    assign OUT[25] = p_0[25] ^ g_8_24;
    assign OUT[26] = p_0[26] ^ g_5_25;
    assign OUT[27] = p_0[27] ^ g_8_26;
    assign OUT[28] = p_0[28] ^ g_5_27;
    assign OUT[29] = p_0[29] ^ g_8_28;
    assign OUT[30] = p_0[30] ^ g_5_29;
    assign OUT[31] = p_0[31] ^ g_8_30;
    assign OUT[32] = p_0[32] ^ g_5_31;
    assign OUT[33] = p_0[33] ^ g_8_32;
    assign OUT[34] = p_0[34] ^ g_6_33;
    assign OUT[35] = p_0[35] ^ g_8_34;
    assign OUT[36] = p_0[36] ^ g_6_35;
    assign OUT[37] = p_0[37] ^ g_8_36;
    assign OUT[38] = p_0[38] ^ g_6_37;
    assign OUT[39] = p_0[39] ^ g_8_38;
    assign OUT[40] = p_0[40] ^ g_6_39;
    assign OUT[41] = p_0[41] ^ g_8_40;
    assign OUT[42] = p_0[42] ^ g_6_41;
    assign OUT[43] = p_0[43] ^ g_8_42;
    assign OUT[44] = p_0[44] ^ g_6_43;
    assign OUT[45] = p_0[45] ^ g_8_44;
    assign OUT[46] = p_0[46] ^ g_6_45;
    assign OUT[47] = p_0[47] ^ g_8_46;
    assign OUT[48] = p_0[48] ^ g_6_47;
    assign OUT[49] = p_0[49] ^ g_8_48;
    assign OUT[50] = p_0[50] ^ g_6_49;
    assign OUT[51] = p_0[51] ^ g_8_50;
    assign OUT[52] = p_0[52] ^ g_6_51;
    assign OUT[53] = p_0[53] ^ g_8_52;
    assign OUT[54] = p_0[54] ^ g_6_53;
    assign OUT[55] = p_0[55] ^ g_8_54;
    assign OUT[56] = p_0[56] ^ g_6_55;
    assign OUT[57] = p_0[57] ^ g_8_56;
    assign OUT[58] = p_0[58] ^ g_6_57;
    assign OUT[59] = p_0[59] ^ g_8_58;
    assign OUT[60] = p_0[60] ^ g_6_59;
    assign OUT[61] = p_0[61] ^ g_8_60;
    assign OUT[62] = p_0[62] ^ g_6_61;
    assign OUT[63] = p_0[63] ^ g_8_62;
    assign OUT[64] = p_0[64] ^ g_6_63;
    assign OUT[65] = p_0[65] ^ g_8_64;
    assign OUT[66] = p_0[66] ^ g_7_65;
    assign OUT[67] = p_0[67] ^ g_8_66;
    assign OUT[68] = p_0[68] ^ g_7_67;
    assign OUT[69] = p_0[69] ^ g_8_68;
    assign OUT[70] = p_0[70] ^ g_7_69;
    assign OUT[71] = p_0[71] ^ g_8_70;
    assign OUT[72] = p_0[72] ^ g_7_71;
    assign OUT[73] = p_0[73] ^ g_8_72;
    assign OUT[74] = p_0[74] ^ g_7_73;
    assign OUT[75] = p_0[75] ^ g_8_74;
    assign OUT[76] = p_0[76] ^ g_7_75;
    assign OUT[77] = p_0[77] ^ g_8_76;
    assign OUT[78] = p_0[78] ^ g_7_77;
    assign OUT[79] = p_0[79] ^ g_8_78;
    assign OUT[80] = p_0[80] ^ g_7_79;
    assign OUT[81] = p_0[81] ^ g_8_80;
    assign OUT[82] = p_0[82] ^ g_7_81;
    assign OUT[83] = p_0[83] ^ g_8_82;
    assign OUT[84] = p_0[84] ^ g_7_83;
    assign OUT[85] = p_0[85] ^ g_8_84;
    assign OUT[86] = p_0[86] ^ g_7_85;
    assign OUT[87] = p_0[87] ^ g_8_86;
    assign OUT[88] = p_0[88] ^ g_7_87;
    assign OUT[89] = p_0[89] ^ g_8_88;
    assign OUT[90] = p_0[90] ^ g_7_89;
    assign OUT[91] = p_0[91] ^ g_8_90;
    assign OUT[92] = p_0[92] ^ g_7_91;
    assign OUT[93] = p_0[93] ^ g_8_92;
    assign OUT[94] = p_0[94] ^ g_7_93;
    assign OUT[95] = p_0[95] ^ g_8_94;
    assign OUT[96] = p_0[96] ^ g_7_95;
    assign OUT[97] = p_0[97] ^ g_8_96;
    assign OUT[98] = p_0[98] ^ g_7_97;
    assign OUT[99] = p_0[99] ^ g_8_98;
    assign OUT[100] = p_0[100] ^ g_7_99;
    assign OUT[101] = p_0[101] ^ g_8_100;
    assign OUT[102] = p_0[102] ^ g_7_101;
    assign OUT[103] = p_0[103] ^ g_8_102;
    assign OUT[104] = p_0[104] ^ g_7_103;
    assign OUT[105] = p_0[105] ^ g_8_104;
    assign OUT[106] = p_0[106] ^ g_7_105;
    assign OUT[107] = p_0[107] ^ g_8_106;
    assign OUT[108] = p_0[108] ^ g_7_107;
    assign OUT[109] = p_0[109] ^ g_8_108;
    assign OUT[110] = p_0[110] ^ g_7_109;
    assign OUT[111] = p_0[111] ^ g_8_110;
    assign OUT[112] = p_0[112] ^ g_7_111;
    assign OUT[113] = p_0[113] ^ g_8_112;
    assign OUT[114] = p_0[114] ^ g_7_113;
    assign OUT[115] = p_0[115] ^ g_8_114;
    assign OUT[116] = p_0[116] ^ g_7_115;
    assign OUT[117] = p_0[117] ^ g_8_116;
    assign OUT[118] = p_0[118] ^ g_7_117;
    assign OUT[119] = p_0[119] ^ g_8_118;
    assign OUT[120] = p_0[120] ^ g_7_119;
    assign OUT[121] = p_0[121] ^ g_8_120;
    assign OUT[122] = p_0[122] ^ g_7_121;
    assign OUT[123] = p_0[123] ^ g_8_122;
    assign OUT[124] = p_0[124] ^ g_7_123;
    assign OUT[125] = p_0[125] ^ g_8_124;
    assign OUT[126] = p_0[126] ^ g_7_125;
    assign OUT[127] = p_0[127] ^ g_8_126;
    assign OUT[128] = g_7_127;
endmodule

