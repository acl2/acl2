
module top ;

// Can't use undefined preprocessor macro
wire w = `foo;

endmodule
