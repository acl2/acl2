

module top ;

  import pack::*; // package doesn't exist

endmodule
