module tricky;
  logic [2:0] foo_t;
endmodule

module top (tricky.foo_t a);

endmodule
