package pack;


endpackage


module top (output topout, input topin);

  import pack::foo;  // does not exist

endmodule
