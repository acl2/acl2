module top () ;

   // oops, forgot to declare foo_t
   //   typedef logic [1:0] foo_t;

   enum foo_t {FOO, BAR} a;

endmodule
