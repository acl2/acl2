// SVEX - Symbolic, Vector-Level Hardware Description Library
// Copyright (C) 2014 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Sol Swords <sswords@centtech.com>

typedef struct packed {
  logic [3:0] a;
  logic [3:0] b;
  logic [3:0] op;
} alu_in;

module sub (input alu_in ain,
	    output logic [3:0] res);

   assign res = ain.op[1] ?
		ain.op[0] ? ain.a + ain.b : ain.a - ain.b :
		ain.op[0] ? ain.a & ain.b : ain.a | ain.b;

endmodule // sub

module spec (input logic [127:0] in,
	     output wire [127:0] out);

   alu_in ain;
   assign ain.a = in[3:0];
   assign ain.b = in[7:4];
   assign ain.op = in[11:8];

   sub subinst (.ain(ain), .res(out[3:0]));

endmodule // spec
