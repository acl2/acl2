// VL Verilog Toolkit
// Copyright (C) 2008-2015 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
//   THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Jared Davis <jared@centtech.com>

// This is just checking some fancy port handling

module m0 #(width = 4, height = 7)
  (output [width-1:0] o,
   input [width-1:0] a,
   input [width-1:0] b);
  assign o = a & b;
endmodule

module m1 (output logic [3:0][4:0] o,  // 4*5 == 20 bits
           input logic [4:0][3:0] a,   // 5*4 == 20 bits
	   input logic [5:0][3:0] b);  // 6*4 == 24 bits
  assign o = a & b;
endmodule

module m2 (output logic [3:0] omega [4:0],
           input logic [3:0] alpha [5:0],
	   input logic [3:0] beta [6:0]);
endmodule

module m3 (output logic [3:0] omega [4],
           input logic [3:0] alpha [5],
	   input logic [3:0] beta [6]);
endmodule
