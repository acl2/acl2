package pack;


endpackage


module top ;

  import pack::foo;  // does not exist

endmodule
