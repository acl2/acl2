module top ;

  sub mysub ();

endmodule


module sub ;



endmodule : oops   // oops, not the right name
