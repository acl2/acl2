module foo ;
  integer a;
  integer b = ++a++;
endmodule
