
module top ();

  function foo (input a) ;
    foo = b;                // oops, b not declared
  endfunction

endmodule

