// VL preprocessor test
// Copyright (C) 2016 Apple, Inc.
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Jared Davis

module spec (input logic [127:0] in,
	     output wire [127:0] out);

   // This is a horrible corner case for the preprocessor.  What does
   // a line continuation expand to?
   //
   //   -- If it expands to nothing or a space or something like that,
   //      then `HORRIBLE should result in `define FOO 1'b1
   //   -- If it expands to a newline, then `HORRIBLE should expand to
   //          `define FOO
   //          1'b1
   //
   // We find that in both NCV and VCS, it seems to behave like a newline.

   `define HORRIBLE \
      `define FOO \
      1'b1

   generate
      if (`HORRIBLE) begin
	 assign out[3:0] = ~in[3:0];
      end
      else begin
	 assign out[3:0] = in[3:0];
      end
   endgenerate

   `ifdef FOO
   assign out[7:4] = ~in[7:4];
   `else
   assign out[7:4] = in[7:4];
   `endif

   assign out[127:8] = '0;

endmodule
