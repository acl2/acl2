/*----------------------------------------------------------------------------
  Copyright (c) 2004 Aoki laboratory. All rights reserved.

  Top module: Multiplier_63_0_6000

  Number system: 2's complement
  Multiplicand length: 64
  Multiplier length: 64
  Partial product generation: PPG with Radix-4 modified Booth recoding
  Partial product accumulation: (7,3) counter tree
  Final stage addition: Carry select adder
----------------------------------------------------------------------------*/

module TCDECON_63_0(TOP, R, I);
  output [62:0] R;
  output [63:63] TOP;
  input [63:0] I;
  assign TOP[63] = I[63];
  assign R[0] = I[0];
  assign R[1] = I[1];
  assign R[2] = I[2];
  assign R[3] = I[3];
  assign R[4] = I[4];
  assign R[5] = I[5];
  assign R[6] = I[6];
  assign R[7] = I[7];
  assign R[8] = I[8];
  assign R[9] = I[9];
  assign R[10] = I[10];
  assign R[11] = I[11];
  assign R[12] = I[12];
  assign R[13] = I[13];
  assign R[14] = I[14];
  assign R[15] = I[15];
  assign R[16] = I[16];
  assign R[17] = I[17];
  assign R[18] = I[18];
  assign R[19] = I[19];
  assign R[20] = I[20];
  assign R[21] = I[21];
  assign R[22] = I[22];
  assign R[23] = I[23];
  assign R[24] = I[24];
  assign R[25] = I[25];
  assign R[26] = I[26];
  assign R[27] = I[27];
  assign R[28] = I[28];
  assign R[29] = I[29];
  assign R[30] = I[30];
  assign R[31] = I[31];
  assign R[32] = I[32];
  assign R[33] = I[33];
  assign R[34] = I[34];
  assign R[35] = I[35];
  assign R[36] = I[36];
  assign R[37] = I[37];
  assign R[38] = I[38];
  assign R[39] = I[39];
  assign R[40] = I[40];
  assign R[41] = I[41];
  assign R[42] = I[42];
  assign R[43] = I[43];
  assign R[44] = I[44];
  assign R[45] = I[45];
  assign R[46] = I[46];
  assign R[47] = I[47];
  assign R[48] = I[48];
  assign R[49] = I[49];
  assign R[50] = I[50];
  assign R[51] = I[51];
  assign R[52] = I[52];
  assign R[53] = I[53];
  assign R[54] = I[54];
  assign R[55] = I[55];
  assign R[56] = I[56];
  assign R[57] = I[57];
  assign R[58] = I[58];
  assign R[59] = I[59];
  assign R[60] = I[60];
  assign R[61] = I[61];
  assign R[62] = I[62];
endmodule

module R4BEEL_0_2(O_ds, O_d1, O_d0, I2, I1);
  output O_ds, O_d1, O_d0;
  input I1;
  input I2;
  assign O_d0 = I1;
  assign O_d1 = I2 & ( ~ I1 );
  assign O_ds = I2;
endmodule

module R4BEE_1(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_2(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_3(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_4(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_5(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_6(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_7(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_8(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_9(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_10(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_11(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_12(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_13(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_14(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_15(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_16(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_17(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_18(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_19(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_20(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_21(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_22(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_23(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_24(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_25(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_26(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_27(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_28(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_29(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEE_30(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module R4BEEH_31_3(O_ds, O_d1, O_d0, I2, I1, I0);
  output O_ds, O_d1, O_d0;
  input I0;
  input I1;
  input I2;
  assign O_d0 = I1 ^ I0;
  assign O_d1 = ( I2 ^ I1 ) & ( ~ ( I1 ^ I0 ) );
  assign O_ds = I2;
endmodule

module SD41DDECON_0(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_0(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_0(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_0(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_1(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_2(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_3(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_4(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_5(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_6(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_7(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_8(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_9(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_10(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_11(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_12(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_13(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_14(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_15(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_16(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_17(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_18(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_19(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_20(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_21(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_22(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_23(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_24(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_25(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_26(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_27(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_28(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_29(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_30(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_31(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_32(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_33(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_34(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_35(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_36(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_37(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_38(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_39(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_40(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_41(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_42(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_43(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_44(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_45(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_46(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_47(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_48(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_49(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_50(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_51(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_52(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_53(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_54(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_55(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_56(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_57(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_58(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_59(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_60(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_61(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_62(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_63(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_64(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_0(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_1(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_1(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_1(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_64(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_65(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_66(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_2(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_2(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_2(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_2(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_66(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_67(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_68(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_4(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_3(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_3(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_3(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_68(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_69(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_70(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_6(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_4(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_4(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_4(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_70(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_71(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_72(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_8(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_5(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_5(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_5(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_72(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_73(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_74(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_10(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_6(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_6(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_6(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_74(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_75(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_76(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_12(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_7(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_7(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_7(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_76(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_77(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_78(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_14(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_8(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_8(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_8(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_78(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_79(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_80(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_16(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_9(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_9(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_9(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_80(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_81(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_82(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_18(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_10(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_10(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_10(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_82(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_83(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_84(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_20(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_11(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_11(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_11(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_84(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_85(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_86(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_22(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_12(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_12(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_12(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_86(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_87(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_88(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_24(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_13(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_13(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_13(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_88(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_89(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_90(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_26(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_14(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_14(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_14(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_90(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_91(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_92(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_28(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_15(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_15(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_15(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_92(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_93(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_94(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_30(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_16(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_16(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_16(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_94(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_95(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_96(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_32(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_17(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_17(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_17(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_96(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_97(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_98(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_34(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_18(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_18(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_18(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_98(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_99(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_100(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_36(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_19(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_19(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_19(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_100(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_101(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_102(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_38(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_20(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_20(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_20(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_102(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_103(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_104(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_40(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_21(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_21(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_21(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_104(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_105(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_106(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_42(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_22(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_22(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_22(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_106(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_107(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_108(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_44(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_23(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_23(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_23(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_108(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_109(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_110(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_46(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_24(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_24(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_24(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_110(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_111(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_112(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_48(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_25(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_25(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_25(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_112(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_113(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_114(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_50(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_26(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_26(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_26(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_114(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_115(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_116(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_52(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_27(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_27(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_27(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_116(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_117(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_118(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_54(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_28(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_28(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_28(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_118(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_119(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_120(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_56(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_29(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_29(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_29(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_120(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_121(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_122(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_58(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_30(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_30(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_30(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_122(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_123(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_124(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_60(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module SD41DDECON_31(S, U_d1, U_d0, I_ds, I_d1, I_d0);
  output S;
  output U_d1, U_d0;
  input I_ds, I_d1, I_d0;
  assign S = I_ds;
  assign U_d0 = I_d0;
  assign U_d1 = I_d1;
endmodule

module U4DPPGL_0_31(Po, O, I, U_d1, U_d0);
  output O;
  output Po;
  input I;
  input U_d1, U_d0;
  assign O = I & U_d0;
  assign Po = I & U_d1;
endmodule

module U4DPPG_1_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_2_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_3_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_4_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_5_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_6_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_7_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_8_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_9_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_10_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_11_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_12_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_13_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_14_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_15_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_16_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_17_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_18_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_19_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_20_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_21_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_22_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_23_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_24_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_25_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_26_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_27_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_28_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_29_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_30_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_31_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_32_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_33_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_34_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_35_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_36_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_37_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_38_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_39_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_40_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_41_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_42_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_43_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_44_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_45_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_46_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_47_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_48_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_49_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_50_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_51_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_52_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_53_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_54_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_55_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_56_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_57_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_58_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_59_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_60_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_61_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPG_62_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & U_d1;
endmodule

module U4DPPGH_63_31(Po, O, I, U_d1, U_d0, Pi);
  output O;
  output Po;
  input I;
  input Pi;
  input U_d1, U_d0;
  assign O = ( I & U_d0 ) | Pi;
  assign Po = I & ( U_d1 | U_d0 );
endmodule

module BWCPP_124(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCPP_125(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ I;
endmodule

module BWCNP_126(O, I, S);
  output O;
  input I;
  input S;
  assign O = ( ~ S ) ^ I;
endmodule

module UBBBG_62(O, S);
  output O;
  input S;
  assign O = S;
endmodule

module UBOne_65(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_65(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_32(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_33(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_34(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_35(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_36(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_37(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_38(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_39(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_40(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_41(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_42(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_43(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_44(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_45(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_46(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_47(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_48(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_49(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_50(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_51(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_52(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_53(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_54(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_55(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_56(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_57(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_58(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_59(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_60(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_61(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_62(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_63(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_64(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBOne_67(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_67(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_66(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module UBOne_69(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_69(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_68(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_3_3(O);
  output [3:3] O;
  assign O[3] = 0;
endmodule

module UBOne_71(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_71(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_70(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_5_5(O);
  output [5:5] O;
  assign O[5] = 0;
endmodule

module UBOne_73(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_73(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_72(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_7_7(O);
  output [7:7] O;
  assign O[7] = 0;
endmodule

module UBOne_75(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_75(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_74(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_9_9(O);
  output [9:9] O;
  assign O[9] = 0;
endmodule

module UBOne_77(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_77(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_76(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_11_11(O);
  output [11:11] O;
  assign O[11] = 0;
endmodule

module UBOne_79(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_79(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_78(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_13_13(O);
  output [13:13] O;
  assign O[13] = 0;
endmodule

module UBOne_81(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_81(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_80(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_15_15(O);
  output [15:15] O;
  assign O[15] = 0;
endmodule

module UBOne_83(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_83(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_82(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_17_17(O);
  output [17:17] O;
  assign O[17] = 0;
endmodule

module UBOne_85(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_85(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_84(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_19_19(O);
  output [19:19] O;
  assign O[19] = 0;
endmodule

module UBOne_87(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_87(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_86(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_21_21(O);
  output [21:21] O;
  assign O[21] = 0;
endmodule

module UBOne_89(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_89(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_88(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_23_23(O);
  output [23:23] O;
  assign O[23] = 0;
endmodule

module UBOne_91(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_91(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_90(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_25_25(O);
  output [25:25] O;
  assign O[25] = 0;
endmodule

module UBOne_93(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_93(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_92(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_27_27(O);
  output [27:27] O;
  assign O[27] = 0;
endmodule

module UBOne_95(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_95(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_94(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_29_29(O);
  output [29:29] O;
  assign O[29] = 0;
endmodule

module UBOne_97(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_97(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_96(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_31_31(O);
  output [31:31] O;
  assign O[31] = 0;
endmodule

module UBOne_99(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_99(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_98(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_33_33(O);
  output [33:33] O;
  assign O[33] = 0;
endmodule

module UBOne_101(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_101(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_100(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_35_35(O);
  output [35:35] O;
  assign O[35] = 0;
endmodule

module UBOne_103(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_103(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_102(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_37_37(O);
  output [37:37] O;
  assign O[37] = 0;
endmodule

module UBOne_105(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_105(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_104(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_39_39(O);
  output [39:39] O;
  assign O[39] = 0;
endmodule

module UBOne_107(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_107(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_106(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_41_41(O);
  output [41:41] O;
  assign O[41] = 0;
endmodule

module UBOne_109(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_109(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_108(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_43_43(O);
  output [43:43] O;
  assign O[43] = 0;
endmodule

module UBOne_111(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_111(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_110(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_45_45(O);
  output [45:45] O;
  assign O[45] = 0;
endmodule

module UBOne_113(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_113(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_112(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_47_47(O);
  output [47:47] O;
  assign O[47] = 0;
endmodule

module UBOne_115(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_115(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_114(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_49_49(O);
  output [49:49] O;
  assign O[49] = 0;
endmodule

module UBOne_117(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_117(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_116(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_51_51(O);
  output [51:51] O;
  assign O[51] = 0;
endmodule

module UBOne_119(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_119(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_118(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_53_53(O);
  output [53:53] O;
  assign O[53] = 0;
endmodule

module UBOne_121(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_121(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_120(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_55_55(O);
  output [55:55] O;
  assign O[55] = 0;
endmodule

module UBOne_123(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_123(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_122(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_57_57(O);
  output [57:57] O;
  assign O[57] = 0;
endmodule

module UBOne_125(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_125(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_124(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_59_59(O);
  output [59:59] O;
  assign O[59] = 0;
endmodule

module UB1DCON_126(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_61_61(O);
  output [61:61] O;
  assign O[61] = 0;
endmodule

module UBOne_64(O);
  output O;
  assign O = 1;
endmodule

module UBZero_63_63(O);
  output [63:63] O;
  assign O[63] = 0;
endmodule

module UBHA_28(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB4_3C30(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C31(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C32(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C33(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C34(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C35(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C36(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_36(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB7_3C37(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_37(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C38(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C38(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C39(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C39(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C40(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C40(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C41(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C41(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C42(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C43(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C44(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_44(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB7_3C45(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_45(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C46(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C46(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C47(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C47(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C48(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C48(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C49(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C49(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C50(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C51(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C52(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_52(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB7_3C53(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_53(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C54(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C54(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C55(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C55(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C56(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C56(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C57(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C57(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C58(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C59(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C60(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_60(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB7_3C61(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_61(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C62(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C62(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C63(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C63(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C64(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C64(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C65(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C65(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C66(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_66(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C67(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_67(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C68(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C69(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C69(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C70(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C70(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C71(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C71(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C72(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C72(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C73(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C73(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C74(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_74(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C75(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_75(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C76(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C77(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C77(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C78(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C78(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C79(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C79(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C80(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C80(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C81(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C81(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C82(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_82(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C83(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_83(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C84(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C85(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C85(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C86(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C86(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C87(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C87(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C88(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C88(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C89(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C89(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C90(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_90(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C91(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_91(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C92(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C93(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C94(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C95(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C96(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C97(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_98(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_99(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB4_3C14(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C15(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C16(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C17(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C18(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C19(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C20(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB7_3C21(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C22(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C22(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C23(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C23(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C24(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C24(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C25(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C25(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C26(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C27(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C28(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C29(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C30(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C31(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C32(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C33(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C93(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C94(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C95(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C96(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C97(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C98(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C99(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C100(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C101(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C101(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C102(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C102(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C103(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C103(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C104(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C104(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C105(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C105(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C106(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_106(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C107(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_107(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C108(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C109(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C110(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C111(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C112(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C113(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_114(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_115(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB4_3C6(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C7(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C8(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C9(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C10(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C11(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C12(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C13(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C14(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C15(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C16(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C17(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C109(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C110(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C111(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C112(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C113(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C114(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C115(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C116(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C117(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C118(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C119(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C120(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C121(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_122(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_123(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_30(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_31(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_32(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_33(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_34(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_35(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_36(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_38(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_39(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_40(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_41(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_42(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_43(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_44(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_46(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_47(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_48(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_49(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_50(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_51(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_52(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_54(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_55(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_56(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_57(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_58(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_59(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_60(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_62(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_63(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_64(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_65(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_68(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_69(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_70(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_71(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_72(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_73(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_76(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_77(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_78(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_79(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_80(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_81(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_84(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_85(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_86(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_87(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_88(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_89(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_92(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_93(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_94(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_95(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_96(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_97(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_100(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_101(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_102(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_103(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_104(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_105(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_108(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_109(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_110(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_111(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_112(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_113(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_116(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_117(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_118(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_119(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_120(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_121(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_124(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_125(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_0(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBOne_1(O);
  output O;
  assign O = 1;
endmodule

module UBFA_1(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSlB_1_1(Co, S, X, Y, Ci);
  output Co;
  output [1:1] S;
  input Ci;
  input [1:1] X;
  input [1:1] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [1:1] S_0;
  wire [1:1] S_1;
  assign S[1] = ( S_0[1] & ( ~ Ci ) ) | ( S_1[1] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_1 U0 (Ci_1);
  UBZero_1_1 U1 (Ci_0);
  UBRCB_1_1 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_1_1 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_2(O);
  output O;
  assign O = 1;
endmodule

module UBZero_2_2(O);
  output [2:2] O;
  assign O[2] = 0;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSlB_3_2(Co, S, X, Y, Ci);
  output Co;
  output [3:2] S;
  input Ci;
  input [3:2] X;
  input [3:2] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [3:2] S_0;
  wire [3:2] S_1;
  assign S[2] = ( S_0[2] & ( ~ Ci ) ) | ( S_1[2] & Ci );
  assign S[3] = ( S_0[3] & ( ~ Ci ) ) | ( S_1[3] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_2 U0 (Ci_1);
  UBZero_2_2 U1 (Ci_0);
  UBRCB_3_2 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_3_2 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_4(O);
  output O;
  assign O = 1;
endmodule

module UBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module UBCSlB_6_4(Co, S, X, Y, Ci);
  output Co;
  output [6:4] S;
  input Ci;
  input [6:4] X;
  input [6:4] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [6:4] S_0;
  wire [6:4] S_1;
  assign S[4] = ( S_0[4] & ( ~ Ci ) ) | ( S_1[4] & Ci );
  assign S[5] = ( S_0[5] & ( ~ Ci ) ) | ( S_1[5] & Ci );
  assign S[6] = ( S_0[6] & ( ~ Ci ) ) | ( S_1[6] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_4 U0 (Ci_1);
  UBZero_4_4 U1 (Ci_0);
  UBRCB_6_4 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_6_4 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_7(O);
  output O;
  assign O = 1;
endmodule

module UBCSlB_10_7(Co, S, X, Y, Ci);
  output Co;
  output [10:7] S;
  input Ci;
  input [10:7] X;
  input [10:7] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [10:7] S_0;
  wire [10:7] S_1;
  assign S[7] = ( S_0[7] & ( ~ Ci ) ) | ( S_1[7] & Ci );
  assign S[8] = ( S_0[8] & ( ~ Ci ) ) | ( S_1[8] & Ci );
  assign S[9] = ( S_0[9] & ( ~ Ci ) ) | ( S_1[9] & Ci );
  assign S[10] = ( S_0[10] & ( ~ Ci ) ) | ( S_1[10] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_7 U0 (Ci_1);
  UBZero_7_7 U1 (Ci_0);
  UBRCB_10_7 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_10_7 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_11(O);
  output O;
  assign O = 1;
endmodule

module UBCSlB_15_11(Co, S, X, Y, Ci);
  output Co;
  output [15:11] S;
  input Ci;
  input [15:11] X;
  input [15:11] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [15:11] S_0;
  wire [15:11] S_1;
  assign S[11] = ( S_0[11] & ( ~ Ci ) ) | ( S_1[11] & Ci );
  assign S[12] = ( S_0[12] & ( ~ Ci ) ) | ( S_1[12] & Ci );
  assign S[13] = ( S_0[13] & ( ~ Ci ) ) | ( S_1[13] & Ci );
  assign S[14] = ( S_0[14] & ( ~ Ci ) ) | ( S_1[14] & Ci );
  assign S[15] = ( S_0[15] & ( ~ Ci ) ) | ( S_1[15] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_11 U0 (Ci_1);
  UBZero_11_11 U1 (Ci_0);
  UBRCB_15_11 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_15_11 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_16(O);
  output O;
  assign O = 1;
endmodule

module UBZero_16_16(O);
  output [16:16] O;
  assign O[16] = 0;
endmodule

module UBCSlB_21_16(Co, S, X, Y, Ci);
  output Co;
  output [21:16] S;
  input Ci;
  input [21:16] X;
  input [21:16] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [21:16] S_0;
  wire [21:16] S_1;
  assign S[16] = ( S_0[16] & ( ~ Ci ) ) | ( S_1[16] & Ci );
  assign S[17] = ( S_0[17] & ( ~ Ci ) ) | ( S_1[17] & Ci );
  assign S[18] = ( S_0[18] & ( ~ Ci ) ) | ( S_1[18] & Ci );
  assign S[19] = ( S_0[19] & ( ~ Ci ) ) | ( S_1[19] & Ci );
  assign S[20] = ( S_0[20] & ( ~ Ci ) ) | ( S_1[20] & Ci );
  assign S[21] = ( S_0[21] & ( ~ Ci ) ) | ( S_1[21] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_16 U0 (Ci_1);
  UBZero_16_16 U1 (Ci_0);
  UBRCB_21_16 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_21_16 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_22(O);
  output O;
  assign O = 1;
endmodule

module UBZero_22_22(O);
  output [22:22] O;
  assign O[22] = 0;
endmodule

module UBCSlB_28_22(Co, S, X, Y, Ci);
  output Co;
  output [28:22] S;
  input Ci;
  input [28:22] X;
  input [28:22] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [28:22] S_0;
  wire [28:22] S_1;
  assign S[22] = ( S_0[22] & ( ~ Ci ) ) | ( S_1[22] & Ci );
  assign S[23] = ( S_0[23] & ( ~ Ci ) ) | ( S_1[23] & Ci );
  assign S[24] = ( S_0[24] & ( ~ Ci ) ) | ( S_1[24] & Ci );
  assign S[25] = ( S_0[25] & ( ~ Ci ) ) | ( S_1[25] & Ci );
  assign S[26] = ( S_0[26] & ( ~ Ci ) ) | ( S_1[26] & Ci );
  assign S[27] = ( S_0[27] & ( ~ Ci ) ) | ( S_1[27] & Ci );
  assign S[28] = ( S_0[28] & ( ~ Ci ) ) | ( S_1[28] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_22 U0 (Ci_1);
  UBZero_22_22 U1 (Ci_0);
  UBRCB_28_22 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_28_22 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_29(O);
  output O;
  assign O = 1;
endmodule

module UBCSlB_36_29(Co, S, X, Y, Ci);
  output Co;
  output [36:29] S;
  input Ci;
  input [36:29] X;
  input [36:29] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [36:29] S_0;
  wire [36:29] S_1;
  assign S[29] = ( S_0[29] & ( ~ Ci ) ) | ( S_1[29] & Ci );
  assign S[30] = ( S_0[30] & ( ~ Ci ) ) | ( S_1[30] & Ci );
  assign S[31] = ( S_0[31] & ( ~ Ci ) ) | ( S_1[31] & Ci );
  assign S[32] = ( S_0[32] & ( ~ Ci ) ) | ( S_1[32] & Ci );
  assign S[33] = ( S_0[33] & ( ~ Ci ) ) | ( S_1[33] & Ci );
  assign S[34] = ( S_0[34] & ( ~ Ci ) ) | ( S_1[34] & Ci );
  assign S[35] = ( S_0[35] & ( ~ Ci ) ) | ( S_1[35] & Ci );
  assign S[36] = ( S_0[36] & ( ~ Ci ) ) | ( S_1[36] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_29 U0 (Ci_1);
  UBZero_29_29 U1 (Ci_0);
  UBRCB_36_29 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_36_29 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_37(O);
  output O;
  assign O = 1;
endmodule

module UBCSlB_45_37(Co, S, X, Y, Ci);
  output Co;
  output [45:37] S;
  input Ci;
  input [45:37] X;
  input [45:37] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [45:37] S_0;
  wire [45:37] S_1;
  assign S[37] = ( S_0[37] & ( ~ Ci ) ) | ( S_1[37] & Ci );
  assign S[38] = ( S_0[38] & ( ~ Ci ) ) | ( S_1[38] & Ci );
  assign S[39] = ( S_0[39] & ( ~ Ci ) ) | ( S_1[39] & Ci );
  assign S[40] = ( S_0[40] & ( ~ Ci ) ) | ( S_1[40] & Ci );
  assign S[41] = ( S_0[41] & ( ~ Ci ) ) | ( S_1[41] & Ci );
  assign S[42] = ( S_0[42] & ( ~ Ci ) ) | ( S_1[42] & Ci );
  assign S[43] = ( S_0[43] & ( ~ Ci ) ) | ( S_1[43] & Ci );
  assign S[44] = ( S_0[44] & ( ~ Ci ) ) | ( S_1[44] & Ci );
  assign S[45] = ( S_0[45] & ( ~ Ci ) ) | ( S_1[45] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_37 U0 (Ci_1);
  UBZero_37_37 U1 (Ci_0);
  UBRCB_45_37 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_45_37 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_46(O);
  output O;
  assign O = 1;
endmodule

module UBZero_46_46(O);
  output [46:46] O;
  assign O[46] = 0;
endmodule

module UBCSlB_55_46(Co, S, X, Y, Ci);
  output Co;
  output [55:46] S;
  input Ci;
  input [55:46] X;
  input [55:46] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [55:46] S_0;
  wire [55:46] S_1;
  assign S[46] = ( S_0[46] & ( ~ Ci ) ) | ( S_1[46] & Ci );
  assign S[47] = ( S_0[47] & ( ~ Ci ) ) | ( S_1[47] & Ci );
  assign S[48] = ( S_0[48] & ( ~ Ci ) ) | ( S_1[48] & Ci );
  assign S[49] = ( S_0[49] & ( ~ Ci ) ) | ( S_1[49] & Ci );
  assign S[50] = ( S_0[50] & ( ~ Ci ) ) | ( S_1[50] & Ci );
  assign S[51] = ( S_0[51] & ( ~ Ci ) ) | ( S_1[51] & Ci );
  assign S[52] = ( S_0[52] & ( ~ Ci ) ) | ( S_1[52] & Ci );
  assign S[53] = ( S_0[53] & ( ~ Ci ) ) | ( S_1[53] & Ci );
  assign S[54] = ( S_0[54] & ( ~ Ci ) ) | ( S_1[54] & Ci );
  assign S[55] = ( S_0[55] & ( ~ Ci ) ) | ( S_1[55] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_46 U0 (Ci_1);
  UBZero_46_46 U1 (Ci_0);
  UBRCB_55_46 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_55_46 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_56(O);
  output O;
  assign O = 1;
endmodule

module UBZero_56_56(O);
  output [56:56] O;
  assign O[56] = 0;
endmodule

module UBCSlB_66_56(Co, S, X, Y, Ci);
  output Co;
  output [66:56] S;
  input Ci;
  input [66:56] X;
  input [66:56] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [66:56] S_0;
  wire [66:56] S_1;
  assign S[56] = ( S_0[56] & ( ~ Ci ) ) | ( S_1[56] & Ci );
  assign S[57] = ( S_0[57] & ( ~ Ci ) ) | ( S_1[57] & Ci );
  assign S[58] = ( S_0[58] & ( ~ Ci ) ) | ( S_1[58] & Ci );
  assign S[59] = ( S_0[59] & ( ~ Ci ) ) | ( S_1[59] & Ci );
  assign S[60] = ( S_0[60] & ( ~ Ci ) ) | ( S_1[60] & Ci );
  assign S[61] = ( S_0[61] & ( ~ Ci ) ) | ( S_1[61] & Ci );
  assign S[62] = ( S_0[62] & ( ~ Ci ) ) | ( S_1[62] & Ci );
  assign S[63] = ( S_0[63] & ( ~ Ci ) ) | ( S_1[63] & Ci );
  assign S[64] = ( S_0[64] & ( ~ Ci ) ) | ( S_1[64] & Ci );
  assign S[65] = ( S_0[65] & ( ~ Ci ) ) | ( S_1[65] & Ci );
  assign S[66] = ( S_0[66] & ( ~ Ci ) ) | ( S_1[66] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_56 U0 (Ci_1);
  UBZero_56_56 U1 (Ci_0);
  UBRCB_66_56 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_66_56 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_67_67(O);
  output [67:67] O;
  assign O[67] = 0;
endmodule

module UBCSlB_78_67(Co, S, X, Y, Ci);
  output Co;
  output [78:67] S;
  input Ci;
  input [78:67] X;
  input [78:67] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [78:67] S_0;
  wire [78:67] S_1;
  assign S[67] = ( S_0[67] & ( ~ Ci ) ) | ( S_1[67] & Ci );
  assign S[68] = ( S_0[68] & ( ~ Ci ) ) | ( S_1[68] & Ci );
  assign S[69] = ( S_0[69] & ( ~ Ci ) ) | ( S_1[69] & Ci );
  assign S[70] = ( S_0[70] & ( ~ Ci ) ) | ( S_1[70] & Ci );
  assign S[71] = ( S_0[71] & ( ~ Ci ) ) | ( S_1[71] & Ci );
  assign S[72] = ( S_0[72] & ( ~ Ci ) ) | ( S_1[72] & Ci );
  assign S[73] = ( S_0[73] & ( ~ Ci ) ) | ( S_1[73] & Ci );
  assign S[74] = ( S_0[74] & ( ~ Ci ) ) | ( S_1[74] & Ci );
  assign S[75] = ( S_0[75] & ( ~ Ci ) ) | ( S_1[75] & Ci );
  assign S[76] = ( S_0[76] & ( ~ Ci ) ) | ( S_1[76] & Ci );
  assign S[77] = ( S_0[77] & ( ~ Ci ) ) | ( S_1[77] & Ci );
  assign S[78] = ( S_0[78] & ( ~ Ci ) ) | ( S_1[78] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_67 U0 (Ci_1);
  UBZero_67_67 U1 (Ci_0);
  UBRCB_78_67 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_78_67 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_79_79(O);
  output [79:79] O;
  assign O[79] = 0;
endmodule

module UBCSlB_91_79(Co, S, X, Y, Ci);
  output Co;
  output [91:79] S;
  input Ci;
  input [91:79] X;
  input [91:79] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [91:79] S_0;
  wire [91:79] S_1;
  assign S[79] = ( S_0[79] & ( ~ Ci ) ) | ( S_1[79] & Ci );
  assign S[80] = ( S_0[80] & ( ~ Ci ) ) | ( S_1[80] & Ci );
  assign S[81] = ( S_0[81] & ( ~ Ci ) ) | ( S_1[81] & Ci );
  assign S[82] = ( S_0[82] & ( ~ Ci ) ) | ( S_1[82] & Ci );
  assign S[83] = ( S_0[83] & ( ~ Ci ) ) | ( S_1[83] & Ci );
  assign S[84] = ( S_0[84] & ( ~ Ci ) ) | ( S_1[84] & Ci );
  assign S[85] = ( S_0[85] & ( ~ Ci ) ) | ( S_1[85] & Ci );
  assign S[86] = ( S_0[86] & ( ~ Ci ) ) | ( S_1[86] & Ci );
  assign S[87] = ( S_0[87] & ( ~ Ci ) ) | ( S_1[87] & Ci );
  assign S[88] = ( S_0[88] & ( ~ Ci ) ) | ( S_1[88] & Ci );
  assign S[89] = ( S_0[89] & ( ~ Ci ) ) | ( S_1[89] & Ci );
  assign S[90] = ( S_0[90] & ( ~ Ci ) ) | ( S_1[90] & Ci );
  assign S[91] = ( S_0[91] & ( ~ Ci ) ) | ( S_1[91] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_79 U0 (Ci_1);
  UBZero_79_79 U1 (Ci_0);
  UBRCB_91_79 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_91_79 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_92(O);
  output O;
  assign O = 1;
endmodule

module UBZero_92_92(O);
  output [92:92] O;
  assign O[92] = 0;
endmodule

module UBCSlB_105_92(Co, S, X, Y, Ci);
  output Co;
  output [105:92] S;
  input Ci;
  input [105:92] X;
  input [105:92] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [105:92] S_0;
  wire [105:92] S_1;
  assign S[92] = ( S_0[92] & ( ~ Ci ) ) | ( S_1[92] & Ci );
  assign S[93] = ( S_0[93] & ( ~ Ci ) ) | ( S_1[93] & Ci );
  assign S[94] = ( S_0[94] & ( ~ Ci ) ) | ( S_1[94] & Ci );
  assign S[95] = ( S_0[95] & ( ~ Ci ) ) | ( S_1[95] & Ci );
  assign S[96] = ( S_0[96] & ( ~ Ci ) ) | ( S_1[96] & Ci );
  assign S[97] = ( S_0[97] & ( ~ Ci ) ) | ( S_1[97] & Ci );
  assign S[98] = ( S_0[98] & ( ~ Ci ) ) | ( S_1[98] & Ci );
  assign S[99] = ( S_0[99] & ( ~ Ci ) ) | ( S_1[99] & Ci );
  assign S[100] = ( S_0[100] & ( ~ Ci ) ) | ( S_1[100] & Ci );
  assign S[101] = ( S_0[101] & ( ~ Ci ) ) | ( S_1[101] & Ci );
  assign S[102] = ( S_0[102] & ( ~ Ci ) ) | ( S_1[102] & Ci );
  assign S[103] = ( S_0[103] & ( ~ Ci ) ) | ( S_1[103] & Ci );
  assign S[104] = ( S_0[104] & ( ~ Ci ) ) | ( S_1[104] & Ci );
  assign S[105] = ( S_0[105] & ( ~ Ci ) ) | ( S_1[105] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_92 U0 (Ci_1);
  UBZero_92_92 U1 (Ci_0);
  UBRCB_105_92 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_105_92 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_106(O);
  output O;
  assign O = 1;
endmodule

module UBZero_106_106(O);
  output [106:106] O;
  assign O[106] = 0;
endmodule

module UBCSlB_120_106(Co, S, X, Y, Ci);
  output Co;
  output [120:106] S;
  input Ci;
  input [120:106] X;
  input [120:106] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [120:106] S_0;
  wire [120:106] S_1;
  assign S[106] = ( S_0[106] & ( ~ Ci ) ) | ( S_1[106] & Ci );
  assign S[107] = ( S_0[107] & ( ~ Ci ) ) | ( S_1[107] & Ci );
  assign S[108] = ( S_0[108] & ( ~ Ci ) ) | ( S_1[108] & Ci );
  assign S[109] = ( S_0[109] & ( ~ Ci ) ) | ( S_1[109] & Ci );
  assign S[110] = ( S_0[110] & ( ~ Ci ) ) | ( S_1[110] & Ci );
  assign S[111] = ( S_0[111] & ( ~ Ci ) ) | ( S_1[111] & Ci );
  assign S[112] = ( S_0[112] & ( ~ Ci ) ) | ( S_1[112] & Ci );
  assign S[113] = ( S_0[113] & ( ~ Ci ) ) | ( S_1[113] & Ci );
  assign S[114] = ( S_0[114] & ( ~ Ci ) ) | ( S_1[114] & Ci );
  assign S[115] = ( S_0[115] & ( ~ Ci ) ) | ( S_1[115] & Ci );
  assign S[116] = ( S_0[116] & ( ~ Ci ) ) | ( S_1[116] & Ci );
  assign S[117] = ( S_0[117] & ( ~ Ci ) ) | ( S_1[117] & Ci );
  assign S[118] = ( S_0[118] & ( ~ Ci ) ) | ( S_1[118] & Ci );
  assign S[119] = ( S_0[119] & ( ~ Ci ) ) | ( S_1[119] & Ci );
  assign S[120] = ( S_0[120] & ( ~ Ci ) ) | ( S_1[120] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_106 U0 (Ci_1);
  UBZero_106_106 U1 (Ci_0);
  UBRCB_120_106 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_120_106 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_121_121(O);
  output [121:121] O;
  assign O[121] = 0;
endmodule

module UBFA_125(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_126(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSlB_126_121(Co, S, X, Y, Ci);
  output Co;
  output [126:121] S;
  input Ci;
  input [126:121] X;
  input [126:121] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [126:121] S_0;
  wire [126:121] S_1;
  assign S[121] = ( S_0[121] & ( ~ Ci ) ) | ( S_1[121] & Ci );
  assign S[122] = ( S_0[122] & ( ~ Ci ) ) | ( S_1[122] & Ci );
  assign S[123] = ( S_0[123] & ( ~ Ci ) ) | ( S_1[123] & Ci );
  assign S[124] = ( S_0[124] & ( ~ Ci ) ) | ( S_1[124] & Ci );
  assign S[125] = ( S_0[125] & ( ~ Ci ) ) | ( S_1[125] & Ci );
  assign S[126] = ( S_0[126] & ( ~ Ci ) ) | ( S_1[126] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_121 U0 (Ci_1);
  UBZero_121_121 U1 (Ci_0);
  UBRCB_126_121 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_126_121 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBPriCSlA_126_0(S, X, Y, Cin);
  output [127:0] S;
  input Cin;
  input [126:0] X;
  input [126:0] Y;
  wire C0;
  wire C1;
  wire C10;
  wire C11;
  wire C12;
  wire C13;
  wire C14;
  wire C15;
  wire C2;
  wire C3;
  wire C4;
  wire C5;
  wire C6;
  wire C7;
  wire C8;
  wire C9;
  UBRCB_0_0 U0 (C0, S[0], X[0], Y[0], Cin);
  UBCSlB_1_1 U1 (C1, S[1], X[1], Y[1], C0);
  UBCSlB_3_2 U2 (C2, S[3:2], X[3:2], Y[3:2], C1);
  UBCSlB_6_4 U3 (C3, S[6:4], X[6:4], Y[6:4], C2);
  UBCSlB_10_7 U4 (C4, S[10:7], X[10:7], Y[10:7], C3);
  UBCSlB_15_11 U5 (C5, S[15:11], X[15:11], Y[15:11], C4);
  UBCSlB_21_16 U6 (C6, S[21:16], X[21:16], Y[21:16], C5);
  UBCSlB_28_22 U7 (C7, S[28:22], X[28:22], Y[28:22], C6);
  UBCSlB_36_29 U8 (C8, S[36:29], X[36:29], Y[36:29], C7);
  UBCSlB_45_37 U9 (C9, S[45:37], X[45:37], Y[45:37], C8);
  UBCSlB_55_46 U10 (C10, S[55:46], X[55:46], Y[55:46], C9);
  UBCSlB_66_56 U11 (C11, S[66:56], X[66:56], Y[66:56], C10);
  UBCSlB_78_67 U12 (C12, S[78:67], X[78:67], Y[78:67], C11);
  UBCSlB_91_79 U13 (C13, S[91:79], X[91:79], Y[91:79], C12);
  UBCSlB_105_92 U14 (C14, S[105:92], X[105:92], Y[105:92], C13);
  UBCSlB_120_106 U15 (C15, S[120:106], X[120:106], Y[120:106], C14);
  UBCSlB_126_121 U16 (S[127], S[126:121], X[126:121], Y[126:121], C15);
endmodule

module UBZero_0_0(O);
  output [0:0] O;
  assign O[0] = 0;
endmodule

module UBTC1CON127_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_32(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_33(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_34(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_35(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_36(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_37(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_38(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_39(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_40(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_41(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_42(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_43(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_44(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_45(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_46(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_47(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_48(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_49(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_50(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_51(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_52(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_53(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_54(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_55(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_56(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_57(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_58(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_59(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_60(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_61(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_62(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_63(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_64(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_65(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_66(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_67(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_68(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_69(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_70(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_71(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_72(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_73(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_74(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_75(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_76(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_77(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_78(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_79(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_80(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_81(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_82(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_83(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_84(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_85(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_86(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_87(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_88(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_89(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_90(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_91(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_92(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_93(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_94(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_95(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_96(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_97(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_98(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_99(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_100(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_101(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_102(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_103(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_104(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_105(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_106(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_107(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_108(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_109(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_110(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_111(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_112(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_113(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_114(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_115(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_116(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_117(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_118(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_119(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_120(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_121(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_122(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_123(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_124(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_125(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON127_126(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTCTCONV_127_127(O, I);
  output [127:127] O;
  input [127:127] I;
  assign O = ~ I;
endmodule

module Multiplier_63_0_6000(P, IN1, IN2);
  output [127:0] P;
  input [63:0] IN1;
  input [63:0] IN2;
  wire [127:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  assign P[28] = W[28];
  assign P[29] = W[29];
  assign P[30] = W[30];
  assign P[31] = W[31];
  assign P[32] = W[32];
  assign P[33] = W[33];
  assign P[34] = W[34];
  assign P[35] = W[35];
  assign P[36] = W[36];
  assign P[37] = W[37];
  assign P[38] = W[38];
  assign P[39] = W[39];
  assign P[40] = W[40];
  assign P[41] = W[41];
  assign P[42] = W[42];
  assign P[43] = W[43];
  assign P[44] = W[44];
  assign P[45] = W[45];
  assign P[46] = W[46];
  assign P[47] = W[47];
  assign P[48] = W[48];
  assign P[49] = W[49];
  assign P[50] = W[50];
  assign P[51] = W[51];
  assign P[52] = W[52];
  assign P[53] = W[53];
  assign P[54] = W[54];
  assign P[55] = W[55];
  assign P[56] = W[56];
  assign P[57] = W[57];
  assign P[58] = W[58];
  assign P[59] = W[59];
  assign P[60] = W[60];
  assign P[61] = W[61];
  assign P[62] = W[62];
  assign P[63] = W[63];
  assign P[64] = W[64];
  assign P[65] = W[65];
  assign P[66] = W[66];
  assign P[67] = W[67];
  assign P[68] = W[68];
  assign P[69] = W[69];
  assign P[70] = W[70];
  assign P[71] = W[71];
  assign P[72] = W[72];
  assign P[73] = W[73];
  assign P[74] = W[74];
  assign P[75] = W[75];
  assign P[76] = W[76];
  assign P[77] = W[77];
  assign P[78] = W[78];
  assign P[79] = W[79];
  assign P[80] = W[80];
  assign P[81] = W[81];
  assign P[82] = W[82];
  assign P[83] = W[83];
  assign P[84] = W[84];
  assign P[85] = W[85];
  assign P[86] = W[86];
  assign P[87] = W[87];
  assign P[88] = W[88];
  assign P[89] = W[89];
  assign P[90] = W[90];
  assign P[91] = W[91];
  assign P[92] = W[92];
  assign P[93] = W[93];
  assign P[94] = W[94];
  assign P[95] = W[95];
  assign P[96] = W[96];
  assign P[97] = W[97];
  assign P[98] = W[98];
  assign P[99] = W[99];
  assign P[100] = W[100];
  assign P[101] = W[101];
  assign P[102] = W[102];
  assign P[103] = W[103];
  assign P[104] = W[104];
  assign P[105] = W[105];
  assign P[106] = W[106];
  assign P[107] = W[107];
  assign P[108] = W[108];
  assign P[109] = W[109];
  assign P[110] = W[110];
  assign P[111] = W[111];
  assign P[112] = W[112];
  assign P[113] = W[113];
  assign P[114] = W[114];
  assign P[115] = W[115];
  assign P[116] = W[116];
  assign P[117] = W[117];
  assign P[118] = W[118];
  assign P[119] = W[119];
  assign P[120] = W[120];
  assign P[121] = W[121];
  assign P[122] = W[122];
  assign P[123] = W[123];
  assign P[124] = W[124];
  assign P[125] = W[125];
  assign P[126] = W[126];
  assign P[127] = W[127];
  MultTC_R4B_D73_CS000 U0 (W, IN1, IN2);
endmodule

module D7_3CTR_126_0_125000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14);
  output [126:0] S1;
  output [126:0] S2;
  input [126:0] PP0;
  input [125:0] PP1;
  input [107:18] PP10;
  input [105:20] PP11;
  input [103:22] PP12;
  input [101:24] PP13;
  input [100:26] PP14;
  input [123:2] PP2;
  input [121:4] PP3;
  input [119:6] PP4;
  input [117:8] PP5;
  input [115:10] PP6;
  input [113:12] PP7;
  input [111:14] PP8;
  input [109:16] PP9;
  wire [126:0] W0;
  wire [125:0] W1;
  wire [123:2] W2;
  wire [121:4] W3;
  wire [119:6] W4;
  wire [117:8] W5;
  wire [116:10] W6;
  UBHA_12 U0 (W5[13], W6[12], PP0[12], PP1[12]);
  UBFA_13 U1 (W5[14], W6[13], PP0[13], PP1[13], PP2[13]);
  UB4_3C14 U2 (W4[16], W5[15], W6[14], PP0[14], PP1[14], PP2[14], PP3[14]);
  UB4_3C15 U3 (W4[17], W5[16], W6[15], PP0[15], PP1[15], PP2[15], PP3[15]);
  UB6_3C16 U4 (W4[18], W5[17], W6[16], PP0[16], PP1[16], PP2[16], PP3[16], PP4[16], PP5[16]);
  UB6_3C17 U5 (W4[19], W5[18], W6[17], PP0[17], PP1[17], PP2[17], PP3[17], PP4[17], PP5[17]);
  UB7_3C18 U6 (W3[20], W5[19], W6[18], PP0[18], PP1[18], PP2[18], PP3[18], PP4[18], PP5[18], PP6[18]);
  UB7_3C19 U7 (W2[21], W4[20], W6[19], PP0[19], PP1[19], PP2[19], PP3[19], PP4[19], PP5[19], PP6[19]);
  UB7_3C20 U8 (W2[22], W3[21], W5[20], PP0[20], PP1[20], PP2[20], PP3[20], PP4[20], PP5[20], PP6[20]);
  UBHA_20 U9 (W4[21], W6[20], PP7[20], PP8[20]);
  UB7_3C21 U10 (W2[23], W3[22], W5[21], PP0[21], PP1[21], PP2[21], PP3[21], PP4[21], PP5[21], PP6[21]);
  UBFA_21 U11 (W4[22], W6[21], PP7[21], PP8[21], PP9[21]);
  UB7_3C22 U12 (W1[24], W3[23], W5[22], PP0[22], PP1[22], PP2[22], PP3[22], PP4[22], PP5[22], PP6[22]);
  UB4_3C22 U13 (W2[24], W4[23], W6[22], PP7[22], PP8[22], PP9[22], PP10[22]);
  UB7_3C23 U14 (W1[25], W3[24], W5[23], PP0[23], PP1[23], PP2[23], PP3[23], PP4[23], PP5[23], PP6[23]);
  UB4_3C23 U15 (W2[25], W4[24], W6[23], PP7[23], PP8[23], PP9[23], PP10[23]);
  UB7_3C24 U16 (W1[26], W3[25], W5[24], PP0[24], PP1[24], PP2[24], PP3[24], PP4[24], PP5[24], PP6[24]);
  UB6_3C24 U17 (W2[26], W4[25], W6[24], PP7[24], PP8[24], PP9[24], PP10[24], PP11[24], PP12[24]);
  UB7_3C25 U18 (W1[27], W3[26], W5[25], PP0[25], PP1[25], PP2[25], PP3[25], PP4[25], PP5[25], PP6[25]);
  UB6_3C25 U19 (W2[27], W4[26], W6[25], PP7[25], PP8[25], PP9[25], PP10[25], PP11[25], PP12[25]);
  UB7_3C26 U20 (W1[28], W3[27], W5[26], PP0[26], PP1[26], PP2[26], PP3[26], PP4[26], PP5[26], PP6[26]);
  UB7_3C26 U21 (W2[28], W4[27], W6[26], PP7[26], PP8[26], PP9[26], PP10[26], PP11[26], PP12[26], PP13[26]);
  UB7_3C27 U22 (W1[29], W3[28], W5[27], PP0[27], PP1[27], PP2[27], PP3[27], PP4[27], PP5[27], PP6[27]);
  UB7_3C27 U23 (W2[29], W4[28], W6[27], PP7[27], PP8[27], PP9[27], PP10[27], PP11[27], PP12[27], PP13[27]);
  UB7_3C28 U24 (W1[30], W3[29], W5[28], PP0[28], PP1[28], PP2[28], PP3[28], PP4[28], PP5[28], PP6[28]);
  UB7_3C28 U25 (W2[30], W4[29], W6[28], PP7[28], PP8[28], PP9[28], PP10[28], PP11[28], PP12[28], PP13[28]);
  UB7_3C29 U26 (W1[31], W3[30], W5[29], PP0[29], PP1[29], PP2[29], PP3[29], PP4[29], PP5[29], PP6[29]);
  UB7_3C29 U27 (W2[31], W4[30], W6[29], PP7[29], PP8[29], PP9[29], PP10[29], PP11[29], PP12[29], PP13[29]);
  UB7_3C30 U28 (W1[32], W3[31], W5[30], PP0[30], PP1[30], PP2[30], PP3[30], PP4[30], PP5[30], PP6[30]);
  UB7_3C30 U29 (W2[32], W4[31], W6[30], PP7[30], PP8[30], PP9[30], PP10[30], PP11[30], PP12[30], PP13[30]);
  UB7_3C31 U30 (W1[33], W3[32], W5[31], PP0[31], PP1[31], PP2[31], PP3[31], PP4[31], PP5[31], PP6[31]);
  UB7_3C31 U31 (W2[33], W4[32], W6[31], PP7[31], PP8[31], PP9[31], PP10[31], PP11[31], PP12[31], PP13[31]);
  UB7_3C32 U32 (W1[34], W3[33], W5[32], PP0[32], PP1[32], PP2[32], PP3[32], PP4[32], PP5[32], PP6[32]);
  UB7_3C32 U33 (W2[34], W4[33], W6[32], PP7[32], PP8[32], PP9[32], PP10[32], PP11[32], PP12[32], PP13[32]);
  UB7_3C33 U34 (W1[35], W3[34], W5[33], PP0[33], PP1[33], PP2[33], PP3[33], PP4[33], PP5[33], PP6[33]);
  UB7_3C33 U35 (W2[35], W4[34], W6[33], PP7[33], PP8[33], PP9[33], PP10[33], PP11[33], PP12[33], PP13[33]);
  UB7_3C34 U36 (W1[36], W3[35], W5[34], PP0[34], PP1[34], PP2[34], PP3[34], PP4[34], PP5[34], PP6[34]);
  UB7_3C34 U37 (W2[36], W4[35], W6[34], PP7[34], PP8[34], PP9[34], PP10[34], PP11[34], PP12[34], PP13[34]);
  UB7_3C35 U38 (W1[37], W3[36], W5[35], PP0[35], PP1[35], PP2[35], PP3[35], PP4[35], PP5[35], PP6[35]);
  UB7_3C35 U39 (W2[37], W4[36], W6[35], PP7[35], PP8[35], PP9[35], PP10[35], PP11[35], PP12[35], PP13[35]);
  UB7_3C36 U40 (W1[38], W3[37], W5[36], PP0[36], PP1[36], PP2[36], PP3[36], PP4[36], PP5[36], PP6[36]);
  UB7_3C36 U41 (W2[38], W4[37], W6[36], PP7[36], PP8[36], PP9[36], PP10[36], PP11[36], PP12[36], PP13[36]);
  UB7_3C37 U42 (W1[39], W3[38], W5[37], PP0[37], PP1[37], PP2[37], PP3[37], PP4[37], PP5[37], PP6[37]);
  UB7_3C37 U43 (W2[39], W4[38], W6[37], PP7[37], PP8[37], PP9[37], PP10[37], PP11[37], PP12[37], PP13[37]);
  UB7_3C38 U44 (W1[40], W3[39], W5[38], PP0[38], PP1[38], PP2[38], PP3[38], PP4[38], PP5[38], PP6[38]);
  UB7_3C38 U45 (W2[40], W4[39], W6[38], PP7[38], PP8[38], PP9[38], PP10[38], PP11[38], PP12[38], PP13[38]);
  UB7_3C39 U46 (W1[41], W3[40], W5[39], PP0[39], PP1[39], PP2[39], PP3[39], PP4[39], PP5[39], PP6[39]);
  UB7_3C39 U47 (W2[41], W4[40], W6[39], PP7[39], PP8[39], PP9[39], PP10[39], PP11[39], PP12[39], PP13[39]);
  UB7_3C40 U48 (W1[42], W3[41], W5[40], PP0[40], PP1[40], PP2[40], PP3[40], PP4[40], PP5[40], PP6[40]);
  UB7_3C40 U49 (W2[42], W4[41], W6[40], PP7[40], PP8[40], PP9[40], PP10[40], PP11[40], PP12[40], PP13[40]);
  UB7_3C41 U50 (W1[43], W3[42], W5[41], PP0[41], PP1[41], PP2[41], PP3[41], PP4[41], PP5[41], PP6[41]);
  UB7_3C41 U51 (W2[43], W4[42], W6[41], PP7[41], PP8[41], PP9[41], PP10[41], PP11[41], PP12[41], PP13[41]);
  UB7_3C42 U52 (W1[44], W3[43], W5[42], PP0[42], PP1[42], PP2[42], PP3[42], PP4[42], PP5[42], PP6[42]);
  UB7_3C42 U53 (W2[44], W4[43], W6[42], PP7[42], PP8[42], PP9[42], PP10[42], PP11[42], PP12[42], PP13[42]);
  UB7_3C43 U54 (W1[45], W3[44], W5[43], PP0[43], PP1[43], PP2[43], PP3[43], PP4[43], PP5[43], PP6[43]);
  UB7_3C43 U55 (W2[45], W4[44], W6[43], PP7[43], PP8[43], PP9[43], PP10[43], PP11[43], PP12[43], PP13[43]);
  UB7_3C44 U56 (W1[46], W3[45], W5[44], PP0[44], PP1[44], PP2[44], PP3[44], PP4[44], PP5[44], PP6[44]);
  UB7_3C44 U57 (W2[46], W4[45], W6[44], PP7[44], PP8[44], PP9[44], PP10[44], PP11[44], PP12[44], PP13[44]);
  UB7_3C45 U58 (W1[47], W3[46], W5[45], PP0[45], PP1[45], PP2[45], PP3[45], PP4[45], PP5[45], PP6[45]);
  UB7_3C45 U59 (W2[47], W4[46], W6[45], PP7[45], PP8[45], PP9[45], PP10[45], PP11[45], PP12[45], PP13[45]);
  UB7_3C46 U60 (W1[48], W3[47], W5[46], PP0[46], PP1[46], PP2[46], PP3[46], PP4[46], PP5[46], PP6[46]);
  UB7_3C46 U61 (W2[48], W4[47], W6[46], PP7[46], PP8[46], PP9[46], PP10[46], PP11[46], PP12[46], PP13[46]);
  UB7_3C47 U62 (W1[49], W3[48], W5[47], PP0[47], PP1[47], PP2[47], PP3[47], PP4[47], PP5[47], PP6[47]);
  UB7_3C47 U63 (W2[49], W4[48], W6[47], PP7[47], PP8[47], PP9[47], PP10[47], PP11[47], PP12[47], PP13[47]);
  UB7_3C48 U64 (W1[50], W3[49], W5[48], PP0[48], PP1[48], PP2[48], PP3[48], PP4[48], PP5[48], PP6[48]);
  UB7_3C48 U65 (W2[50], W4[49], W6[48], PP7[48], PP8[48], PP9[48], PP10[48], PP11[48], PP12[48], PP13[48]);
  UB7_3C49 U66 (W1[51], W3[50], W5[49], PP0[49], PP1[49], PP2[49], PP3[49], PP4[49], PP5[49], PP6[49]);
  UB7_3C49 U67 (W2[51], W4[50], W6[49], PP7[49], PP8[49], PP9[49], PP10[49], PP11[49], PP12[49], PP13[49]);
  UB7_3C50 U68 (W1[52], W3[51], W5[50], PP0[50], PP1[50], PP2[50], PP3[50], PP4[50], PP5[50], PP6[50]);
  UB7_3C50 U69 (W2[52], W4[51], W6[50], PP7[50], PP8[50], PP9[50], PP10[50], PP11[50], PP12[50], PP13[50]);
  UB7_3C51 U70 (W1[53], W3[52], W5[51], PP0[51], PP1[51], PP2[51], PP3[51], PP4[51], PP5[51], PP6[51]);
  UB7_3C51 U71 (W2[53], W4[52], W6[51], PP7[51], PP8[51], PP9[51], PP10[51], PP11[51], PP12[51], PP13[51]);
  UB7_3C52 U72 (W1[54], W3[53], W5[52], PP0[52], PP1[52], PP2[52], PP3[52], PP4[52], PP5[52], PP6[52]);
  UB7_3C52 U73 (W2[54], W4[53], W6[52], PP7[52], PP8[52], PP9[52], PP10[52], PP11[52], PP12[52], PP13[52]);
  UB7_3C53 U74 (W1[55], W3[54], W5[53], PP0[53], PP1[53], PP2[53], PP3[53], PP4[53], PP5[53], PP6[53]);
  UB7_3C53 U75 (W2[55], W4[54], W6[53], PP7[53], PP8[53], PP9[53], PP10[53], PP11[53], PP12[53], PP13[53]);
  UB7_3C54 U76 (W1[56], W3[55], W5[54], PP0[54], PP1[54], PP2[54], PP3[54], PP4[54], PP5[54], PP6[54]);
  UB7_3C54 U77 (W2[56], W4[55], W6[54], PP7[54], PP8[54], PP9[54], PP10[54], PP11[54], PP12[54], PP13[54]);
  UB7_3C55 U78 (W1[57], W3[56], W5[55], PP0[55], PP1[55], PP2[55], PP3[55], PP4[55], PP5[55], PP6[55]);
  UB7_3C55 U79 (W2[57], W4[56], W6[55], PP7[55], PP8[55], PP9[55], PP10[55], PP11[55], PP12[55], PP13[55]);
  UB7_3C56 U80 (W1[58], W3[57], W5[56], PP0[56], PP1[56], PP2[56], PP3[56], PP4[56], PP5[56], PP6[56]);
  UB7_3C56 U81 (W2[58], W4[57], W6[56], PP7[56], PP8[56], PP9[56], PP10[56], PP11[56], PP12[56], PP13[56]);
  UB7_3C57 U82 (W1[59], W3[58], W5[57], PP0[57], PP1[57], PP2[57], PP3[57], PP4[57], PP5[57], PP6[57]);
  UB7_3C57 U83 (W2[59], W4[58], W6[57], PP7[57], PP8[57], PP9[57], PP10[57], PP11[57], PP12[57], PP13[57]);
  UB7_3C58 U84 (W1[60], W3[59], W5[58], PP0[58], PP1[58], PP2[58], PP3[58], PP4[58], PP5[58], PP6[58]);
  UB7_3C58 U85 (W2[60], W4[59], W6[58], PP7[58], PP8[58], PP9[58], PP10[58], PP11[58], PP12[58], PP13[58]);
  UB7_3C59 U86 (W1[61], W3[60], W5[59], PP0[59], PP1[59], PP2[59], PP3[59], PP4[59], PP5[59], PP6[59]);
  UB7_3C59 U87 (W2[61], W4[60], W6[59], PP7[59], PP8[59], PP9[59], PP10[59], PP11[59], PP12[59], PP13[59]);
  UB7_3C60 U88 (W1[62], W3[61], W5[60], PP0[60], PP1[60], PP2[60], PP3[60], PP4[60], PP5[60], PP6[60]);
  UB7_3C60 U89 (W2[62], W4[61], W6[60], PP7[60], PP8[60], PP9[60], PP10[60], PP11[60], PP12[60], PP13[60]);
  UB7_3C61 U90 (W1[63], W3[62], W5[61], PP0[61], PP1[61], PP2[61], PP3[61], PP4[61], PP5[61], PP6[61]);
  UB7_3C61 U91 (W2[63], W4[62], W6[61], PP7[61], PP8[61], PP9[61], PP10[61], PP11[61], PP12[61], PP13[61]);
  UB7_3C62 U92 (W1[64], W3[63], W5[62], PP0[62], PP1[62], PP2[62], PP3[62], PP4[62], PP5[62], PP6[62]);
  UB7_3C62 U93 (W2[64], W4[63], W6[62], PP7[62], PP8[62], PP9[62], PP10[62], PP11[62], PP12[62], PP13[62]);
  UB7_3C63 U94 (W1[65], W3[64], W5[63], PP0[63], PP1[63], PP2[63], PP3[63], PP4[63], PP5[63], PP6[63]);
  UB7_3C63 U95 (W2[65], W4[64], W6[63], PP7[63], PP8[63], PP9[63], PP10[63], PP11[63], PP12[63], PP13[63]);
  UB7_3C64 U96 (W1[66], W3[65], W5[64], PP0[64], PP1[64], PP2[64], PP3[64], PP4[64], PP5[64], PP6[64]);
  UB7_3C64 U97 (W2[66], W4[65], W6[64], PP7[64], PP8[64], PP9[64], PP10[64], PP11[64], PP12[64], PP13[64]);
  UB7_3C65 U98 (W1[67], W3[66], W5[65], PP0[65], PP1[65], PP2[65], PP3[65], PP4[65], PP5[65], PP6[65]);
  UB7_3C65 U99 (W2[67], W4[66], W6[65], PP7[65], PP8[65], PP9[65], PP10[65], PP11[65], PP12[65], PP13[65]);
  UB7_3C66 U100 (W1[68], W3[67], W5[66], PP0[66], PP1[66], PP2[66], PP3[66], PP4[66], PP5[66], PP6[66]);
  UB7_3C66 U101 (W2[68], W4[67], W6[66], PP7[66], PP8[66], PP9[66], PP10[66], PP11[66], PP12[66], PP13[66]);
  UB7_3C67 U102 (W1[69], W3[68], W5[67], PP0[67], PP1[67], PP2[67], PP3[67], PP4[67], PP5[67], PP6[67]);
  UB7_3C67 U103 (W2[69], W4[68], W6[67], PP7[67], PP8[67], PP9[67], PP10[67], PP11[67], PP12[67], PP13[67]);
  UB7_3C68 U104 (W1[70], W3[69], W5[68], PP0[68], PP1[68], PP2[68], PP3[68], PP4[68], PP5[68], PP6[68]);
  UB7_3C68 U105 (W2[70], W4[69], W6[68], PP7[68], PP8[68], PP9[68], PP10[68], PP11[68], PP12[68], PP13[68]);
  UB7_3C69 U106 (W1[71], W3[70], W5[69], PP0[69], PP1[69], PP2[69], PP3[69], PP4[69], PP5[69], PP6[69]);
  UB7_3C69 U107 (W2[71], W4[70], W6[69], PP7[69], PP8[69], PP9[69], PP10[69], PP11[69], PP12[69], PP13[69]);
  UB7_3C70 U108 (W1[72], W3[71], W5[70], PP0[70], PP1[70], PP2[70], PP3[70], PP4[70], PP5[70], PP6[70]);
  UB7_3C70 U109 (W2[72], W4[71], W6[70], PP7[70], PP8[70], PP9[70], PP10[70], PP11[70], PP12[70], PP13[70]);
  UB7_3C71 U110 (W1[73], W3[72], W5[71], PP0[71], PP1[71], PP2[71], PP3[71], PP4[71], PP5[71], PP6[71]);
  UB7_3C71 U111 (W2[73], W4[72], W6[71], PP7[71], PP8[71], PP9[71], PP10[71], PP11[71], PP12[71], PP13[71]);
  UB7_3C72 U112 (W1[74], W3[73], W5[72], PP0[72], PP1[72], PP2[72], PP3[72], PP4[72], PP5[72], PP6[72]);
  UB7_3C72 U113 (W2[74], W4[73], W6[72], PP7[72], PP8[72], PP9[72], PP10[72], PP11[72], PP12[72], PP13[72]);
  UB7_3C73 U114 (W1[75], W3[74], W5[73], PP0[73], PP1[73], PP2[73], PP3[73], PP4[73], PP5[73], PP6[73]);
  UB7_3C73 U115 (W2[75], W4[74], W6[73], PP7[73], PP8[73], PP9[73], PP10[73], PP11[73], PP12[73], PP13[73]);
  UB7_3C74 U116 (W1[76], W3[75], W5[74], PP0[74], PP1[74], PP2[74], PP3[74], PP4[74], PP5[74], PP6[74]);
  UB7_3C74 U117 (W2[76], W4[75], W6[74], PP7[74], PP8[74], PP9[74], PP10[74], PP11[74], PP12[74], PP13[74]);
  UB7_3C75 U118 (W1[77], W3[76], W5[75], PP0[75], PP1[75], PP2[75], PP3[75], PP4[75], PP5[75], PP6[75]);
  UB7_3C75 U119 (W2[77], W4[76], W6[75], PP7[75], PP8[75], PP9[75], PP10[75], PP11[75], PP12[75], PP13[75]);
  UB7_3C76 U120 (W1[78], W3[77], W5[76], PP0[76], PP1[76], PP2[76], PP3[76], PP4[76], PP5[76], PP6[76]);
  UB7_3C76 U121 (W2[78], W4[77], W6[76], PP7[76], PP8[76], PP9[76], PP10[76], PP11[76], PP12[76], PP13[76]);
  UB7_3C77 U122 (W1[79], W3[78], W5[77], PP0[77], PP1[77], PP2[77], PP3[77], PP4[77], PP5[77], PP6[77]);
  UB7_3C77 U123 (W2[79], W4[78], W6[77], PP7[77], PP8[77], PP9[77], PP10[77], PP11[77], PP12[77], PP13[77]);
  UB7_3C78 U124 (W1[80], W3[79], W5[78], PP0[78], PP1[78], PP2[78], PP3[78], PP4[78], PP5[78], PP6[78]);
  UB7_3C78 U125 (W2[80], W4[79], W6[78], PP7[78], PP8[78], PP9[78], PP10[78], PP11[78], PP12[78], PP13[78]);
  UB7_3C79 U126 (W1[81], W3[80], W5[79], PP0[79], PP1[79], PP2[79], PP3[79], PP4[79], PP5[79], PP6[79]);
  UB7_3C79 U127 (W2[81], W4[80], W6[79], PP7[79], PP8[79], PP9[79], PP10[79], PP11[79], PP12[79], PP13[79]);
  UB7_3C80 U128 (W1[82], W3[81], W5[80], PP0[80], PP1[80], PP2[80], PP3[80], PP4[80], PP5[80], PP6[80]);
  UB7_3C80 U129 (W2[82], W4[81], W6[80], PP7[80], PP8[80], PP9[80], PP10[80], PP11[80], PP12[80], PP13[80]);
  UB7_3C81 U130 (W1[83], W3[82], W5[81], PP0[81], PP1[81], PP2[81], PP3[81], PP4[81], PP5[81], PP6[81]);
  UB7_3C81 U131 (W2[83], W4[82], W6[81], PP7[81], PP8[81], PP9[81], PP10[81], PP11[81], PP12[81], PP13[81]);
  UB7_3C82 U132 (W1[84], W3[83], W5[82], PP0[82], PP1[82], PP2[82], PP3[82], PP4[82], PP5[82], PP6[82]);
  UB7_3C82 U133 (W2[84], W4[83], W6[82], PP7[82], PP8[82], PP9[82], PP10[82], PP11[82], PP12[82], PP13[82]);
  UB7_3C83 U134 (W1[85], W3[84], W5[83], PP0[83], PP1[83], PP2[83], PP3[83], PP4[83], PP5[83], PP6[83]);
  UB7_3C83 U135 (W2[85], W4[84], W6[83], PP7[83], PP8[83], PP9[83], PP10[83], PP11[83], PP12[83], PP13[83]);
  UB7_3C84 U136 (W1[86], W3[85], W5[84], PP0[84], PP1[84], PP2[84], PP3[84], PP4[84], PP5[84], PP6[84]);
  UB7_3C84 U137 (W2[86], W4[85], W6[84], PP7[84], PP8[84], PP9[84], PP10[84], PP11[84], PP12[84], PP13[84]);
  UB7_3C85 U138 (W1[87], W3[86], W5[85], PP0[85], PP1[85], PP2[85], PP3[85], PP4[85], PP5[85], PP6[85]);
  UB7_3C85 U139 (W2[87], W4[86], W6[85], PP7[85], PP8[85], PP9[85], PP10[85], PP11[85], PP12[85], PP13[85]);
  UB7_3C86 U140 (W1[88], W3[87], W5[86], PP0[86], PP1[86], PP2[86], PP3[86], PP4[86], PP5[86], PP6[86]);
  UB7_3C86 U141 (W2[88], W4[87], W6[86], PP7[86], PP8[86], PP9[86], PP10[86], PP11[86], PP12[86], PP13[86]);
  UB7_3C87 U142 (W1[89], W3[88], W5[87], PP0[87], PP1[87], PP2[87], PP3[87], PP4[87], PP5[87], PP6[87]);
  UB7_3C87 U143 (W2[89], W4[88], W6[87], PP7[87], PP8[87], PP9[87], PP10[87], PP11[87], PP12[87], PP13[87]);
  UB7_3C88 U144 (W1[90], W3[89], W5[88], PP0[88], PP1[88], PP2[88], PP3[88], PP4[88], PP5[88], PP6[88]);
  UB7_3C88 U145 (W2[90], W4[89], W6[88], PP7[88], PP8[88], PP9[88], PP10[88], PP11[88], PP12[88], PP13[88]);
  UB7_3C89 U146 (W1[91], W3[90], W5[89], PP0[89], PP1[89], PP2[89], PP3[89], PP4[89], PP5[89], PP6[89]);
  UB7_3C89 U147 (W2[91], W4[90], W6[89], PP7[89], PP8[89], PP9[89], PP10[89], PP11[89], PP12[89], PP13[89]);
  UB7_3C90 U148 (W1[92], W3[91], W5[90], PP0[90], PP1[90], PP2[90], PP3[90], PP4[90], PP5[90], PP6[90]);
  UB7_3C90 U149 (W2[92], W4[91], W6[90], PP7[90], PP8[90], PP9[90], PP10[90], PP11[90], PP12[90], PP13[90]);
  UB7_3C91 U150 (W1[93], W3[92], W5[91], PP0[91], PP1[91], PP2[91], PP3[91], PP4[91], PP5[91], PP6[91]);
  UB7_3C91 U151 (W2[93], W4[92], W6[91], PP7[91], PP8[91], PP9[91], PP10[91], PP11[91], PP12[91], PP13[91]);
  UB7_3C92 U152 (W1[94], W3[93], W5[92], PP0[92], PP1[92], PP2[92], PP3[92], PP4[92], PP5[92], PP6[92]);
  UB7_3C92 U153 (W2[94], W4[93], W6[92], PP7[92], PP8[92], PP9[92], PP10[92], PP11[92], PP12[92], PP13[92]);
  UB7_3C93 U154 (W1[95], W3[94], W5[93], PP0[93], PP1[93], PP2[93], PP3[93], PP4[93], PP5[93], PP6[93]);
  UB7_3C93 U155 (W2[95], W4[94], W6[93], PP7[93], PP8[93], PP9[93], PP10[93], PP11[93], PP12[93], PP13[93]);
  UB7_3C94 U156 (W1[96], W3[95], W5[94], PP0[94], PP1[94], PP2[94], PP3[94], PP4[94], PP5[94], PP6[94]);
  UB7_3C94 U157 (W2[96], W4[95], W6[94], PP7[94], PP8[94], PP9[94], PP10[94], PP11[94], PP12[94], PP13[94]);
  UB7_3C95 U158 (W1[97], W3[96], W5[95], PP0[95], PP1[95], PP2[95], PP3[95], PP4[95], PP5[95], PP6[95]);
  UB7_3C95 U159 (W2[97], W4[96], W6[95], PP7[95], PP8[95], PP9[95], PP10[95], PP11[95], PP12[95], PP13[95]);
  UB7_3C96 U160 (W1[98], W3[97], W5[96], PP0[96], PP1[96], PP2[96], PP3[96], PP4[96], PP5[96], PP6[96]);
  UB7_3C96 U161 (W2[98], W4[97], W6[96], PP7[96], PP8[96], PP9[96], PP10[96], PP11[96], PP12[96], PP13[96]);
  UB7_3C97 U162 (W1[99], W3[98], W5[97], PP0[97], PP1[97], PP2[97], PP3[97], PP4[97], PP5[97], PP6[97]);
  UB7_3C97 U163 (W2[99], W4[98], W6[97], PP7[97], PP8[97], PP9[97], PP10[97], PP11[97], PP12[97], PP13[97]);
  UB7_3C98 U164 (W1[100], W3[99], W5[98], PP0[98], PP1[98], PP2[98], PP3[98], PP4[98], PP5[98], PP6[98]);
  UB7_3C98 U165 (W2[100], W4[99], W6[98], PP7[98], PP8[98], PP9[98], PP10[98], PP11[98], PP12[98], PP13[98]);
  UB7_3C99 U166 (W1[101], W3[100], W5[99], PP0[99], PP1[99], PP2[99], PP3[99], PP4[99], PP5[99], PP6[99]);
  UB7_3C99 U167 (W2[101], W4[100], W6[99], PP7[99], PP8[99], PP9[99], PP10[99], PP11[99], PP12[99], PP13[99]);
  UB7_3C100 U168 (W1[102], W3[101], W5[100], PP0[100], PP1[100], PP2[100], PP3[100], PP4[100], PP5[100], PP6[100]);
  UB7_3C100 U169 (W2[102], W4[101], W6[100], PP7[100], PP8[100], PP9[100], PP10[100], PP11[100], PP12[100], PP13[100]);
  UB7_3C101 U170 (W1[103], W3[102], W5[101], PP0[101], PP1[101], PP2[101], PP3[101], PP4[101], PP5[101], PP6[101]);
  UB6_3C101 U171 (W2[103], W4[102], W6[101], PP7[101], PP8[101], PP9[101], PP10[101], PP11[101], PP12[101]);
  UB7_3C102 U172 (W1[104], W3[103], W5[102], PP0[102], PP1[102], PP2[102], PP3[102], PP4[102], PP5[102], PP6[102]);
  UB5_3C102 U173 (W2[104], W4[103], W6[102], PP7[102], PP8[102], PP9[102], PP10[102], PP11[102]);
  UB7_3C103 U174 (W1[105], W3[104], W5[103], PP0[103], PP1[103], PP2[103], PP3[103], PP4[103], PP5[103], PP6[103]);
  UB5_3C103 U175 (W2[105], W4[104], W6[103], PP7[103], PP8[103], PP9[103], PP10[103], PP11[103]);
  UB7_3C104 U176 (W1[106], W3[105], W5[104], PP0[104], PP1[104], PP2[104], PP3[104], PP4[104], PP5[104], PP6[104]);
  UB4_3C104 U177 (W2[106], W4[105], W6[104], PP7[104], PP8[104], PP9[104], PP10[104]);
  UB7_3C105 U178 (W1[107], W3[106], W5[105], PP0[105], PP1[105], PP2[105], PP3[105], PP4[105], PP5[105], PP6[105]);
  UB4_3C105 U179 (W2[107], W4[106], W6[105], PP7[105], PP8[105], PP9[105], PP10[105]);
  UB7_3C106 U180 (W3[108], W3[107], W5[106], PP0[106], PP1[106], PP2[106], PP3[106], PP4[106], PP5[106], PP6[106]);
  UBFA_106 U181 (W4[107], W6[106], PP7[106], PP8[106], PP9[106]);
  UB7_3C107 U182 (W4[109], W4[108], W5[107], PP0[107], PP1[107], PP2[107], PP3[107], PP4[107], PP5[107], PP6[107]);
  UBFA_107 U183 (W5[108], W6[107], PP7[107], PP8[107], PP9[107]);
  UB7_3C108 U184 (W4[110], W5[109], W6[108], PP0[108], PP1[108], PP2[108], PP3[108], PP4[108], PP5[108], PP6[108]);
  UB6_3C109 U185 (W4[111], W5[110], W6[109], PP0[109], PP1[109], PP2[109], PP3[109], PP4[109], PP5[109]);
  UB5_3C110 U186 (W4[112], W5[111], W6[110], PP0[110], PP1[110], PP2[110], PP3[110], PP4[110]);
  UB5_3C111 U187 (W4[113], W5[112], W6[111], PP0[111], PP1[111], PP2[111], PP3[111], PP4[111]);
  UB4_3C112 U188 (W4[114], W5[113], W6[112], PP0[112], PP1[112], PP2[112], PP3[112]);
  UB4_3C113 U189 (W4[115], W5[114], W6[113], PP0[113], PP1[113], PP2[113], PP3[113]);
  UBFA_114 U190 (W5[115], W6[114], PP0[114], PP1[114], PP2[114]);
  UBFA_115 U191 (W6[116], W6[115], PP0[115], PP1[115], PP2[115]);
  UBCON_11_0 U192 (W0[11:0], PP0[11:0]);
  UB1DCON_12 U193 (W0[12], PP2[12]);
  UB1DCON_13 U194 (W0[13], PP3[13]);
  UBCON_15_14 U195 (W0[15:14], PP4[15:14]);
  UBCON_17_16 U196 (W0[17:16], PP6[17:16]);
  UBCON_19_18 U197 (W0[19:18], PP7[19:18]);
  UB1DCON_20 U198 (W0[20], PP9[20]);
  UB1DCON_21 U199 (W0[21], PP10[21]);
  UBCON_23_22 U200 (W0[23:22], PP11[23:22]);
  UBCON_25_24 U201 (W0[25:24], PP13[25:24]);
  UBCON_100_26 U202 (W0[100:26], PP14[100:26]);
  UB1DCON_101 U203 (W0[101], PP13[101]);
  UBCON_103_102 U204 (W0[103:102], PP12[103:102]);
  UBCON_105_104 U205 (W0[105:104], PP11[105:104]);
  UBCON_107_106 U206 (W0[107:106], PP10[107:106]);
  UB1DCON_108 U207 (W0[108], PP7[108]);
  UB1DCON_109 U208 (W0[109], PP6[109]);
  UBCON_111_110 U209 (W0[111:110], PP5[111:110]);
  UBCON_113_112 U210 (W0[113:112], PP4[113:112]);
  UBCON_115_114 U211 (W0[115:114], PP3[115:114]);
  UBCON_126_116 U212 (W0[126:116], PP0[126:116]);
  UBCON_11_0 U213 (W1[11:0], PP1[11:0]);
  UB1DCON_12 U214 (W1[12], PP3[12]);
  UB1DCON_13 U215 (W1[13], PP4[13]);
  UBCON_15_14 U216 (W1[15:14], PP5[15:14]);
  UBCON_17_16 U217 (W1[17:16], PP7[17:16]);
  UBCON_19_18 U218 (W1[19:18], PP8[19:18]);
  UB1DCON_20 U219 (W1[20], PP10[20]);
  UB1DCON_21 U220 (W1[21], PP11[21]);
  UBCON_23_22 U221 (W1[23:22], PP12[23:22]);
  UB1DCON_108 U222 (W1[108], PP8[108]);
  UB1DCON_109 U223 (W1[109], PP7[109]);
  UBCON_111_110 U224 (W1[111:110], PP6[111:110]);
  UBCON_113_112 U225 (W1[113:112], PP5[113:112]);
  UBCON_115_114 U226 (W1[115:114], PP4[115:114]);
  UBCON_125_116 U227 (W1[125:116], PP1[125:116]);
  UBCON_11_2 U228 (W2[11:2], PP2[11:2]);
  UB1DCON_12 U229 (W2[12], PP4[12]);
  UB1DCON_13 U230 (W2[13], PP5[13]);
  UBCON_15_14 U231 (W2[15:14], PP6[15:14]);
  UBCON_17_16 U232 (W2[17:16], PP8[17:16]);
  UBCON_19_18 U233 (W2[19:18], PP9[19:18]);
  UB1DCON_20 U234 (W2[20], PP11[20]);
  UB1DCON_108 U235 (W2[108], PP9[108]);
  UB1DCON_109 U236 (W2[109], PP8[109]);
  UBCON_111_110 U237 (W2[111:110], PP7[111:110]);
  UBCON_113_112 U238 (W2[113:112], PP6[113:112]);
  UBCON_115_114 U239 (W2[115:114], PP5[115:114]);
  UBCON_123_116 U240 (W2[123:116], PP2[123:116]);
  UBCON_11_4 U241 (W3[11:4], PP3[11:4]);
  UB1DCON_12 U242 (W3[12], PP5[12]);
  UB1DCON_13 U243 (W3[13], PP6[13]);
  UBCON_15_14 U244 (W3[15:14], PP7[15:14]);
  UBCON_17_16 U245 (W3[17:16], PP9[17:16]);
  UBCON_19_18 U246 (W3[19:18], PP10[19:18]);
  UB1DCON_109 U247 (W3[109], PP9[109]);
  UBCON_111_110 U248 (W3[111:110], PP8[111:110]);
  UBCON_113_112 U249 (W3[113:112], PP7[113:112]);
  UBCON_115_114 U250 (W3[115:114], PP6[115:114]);
  UBCON_121_116 U251 (W3[121:116], PP3[121:116]);
  UBCON_11_6 U252 (W4[11:6], PP4[11:6]);
  UB1DCON_12 U253 (W4[12], PP6[12]);
  UB1DCON_13 U254 (W4[13], PP7[13]);
  UBCON_15_14 U255 (W4[15:14], PP8[15:14]);
  UBCON_119_116 U256 (W4[119:116], PP4[119:116]);
  UBCON_11_8 U257 (W5[11:8], PP5[11:8]);
  UB1DCON_12 U258 (W5[12], PP7[12]);
  UBCON_117_116 U259 (W5[117:116], PP5[117:116]);
  UBCON_11_10 U260 (W6[11:10], PP6[11:10]);
  D7_3CTR_126_0_125001 U261 (S1, S2, W0, W1, W2, W3, W4, W5, W6);
endmodule

module D7_3CTR_126_0_125001 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6);
  output [126:0] S1;
  output [126:0] S2;
  input [126:0] PP0;
  input [125:0] PP1;
  input [123:2] PP2;
  input [121:4] PP3;
  input [119:6] PP4;
  input [117:8] PP5;
  input [116:10] PP6;
  wire [126:0] W0;
  wire [125:0] W1;
  wire [124:2] W2;
  UBHA_4 U0 (W1[5], W2[4], PP0[4], PP1[4]);
  UBFA_5 U1 (W1[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UB4_3C6 U2 (W0[8], W1[7], W2[6], PP0[6], PP1[6], PP2[6], PP3[6]);
  UB4_3C7 U3 (W0[9], W1[8], W2[7], PP0[7], PP1[7], PP2[7], PP3[7]);
  UB6_3C8 U4 (W0[10], W1[9], W2[8], PP0[8], PP1[8], PP2[8], PP3[8], PP4[8], PP5[8]);
  UB6_3C9 U5 (W0[11], W1[10], W2[9], PP0[9], PP1[9], PP2[9], PP3[9], PP4[9], PP5[9]);
  UB7_3C10 U6 (W0[12], W1[11], W2[10], PP0[10], PP1[10], PP2[10], PP3[10], PP4[10], PP5[10], PP6[10]);
  UB7_3C11 U7 (W0[13], W1[12], W2[11], PP0[11], PP1[11], PP2[11], PP3[11], PP4[11], PP5[11], PP6[11]);
  UB7_3C12 U8 (W0[14], W1[13], W2[12], PP0[12], PP1[12], PP2[12], PP3[12], PP4[12], PP5[12], PP6[12]);
  UB7_3C13 U9 (W0[15], W1[14], W2[13], PP0[13], PP1[13], PP2[13], PP3[13], PP4[13], PP5[13], PP6[13]);
  UB7_3C14 U10 (W0[16], W1[15], W2[14], PP0[14], PP1[14], PP2[14], PP3[14], PP4[14], PP5[14], PP6[14]);
  UB7_3C15 U11 (W0[17], W1[16], W2[15], PP0[15], PP1[15], PP2[15], PP3[15], PP4[15], PP5[15], PP6[15]);
  UB7_3C16 U12 (W0[18], W1[17], W2[16], PP0[16], PP1[16], PP2[16], PP3[16], PP4[16], PP5[16], PP6[16]);
  UB7_3C17 U13 (W0[19], W1[18], W2[17], PP0[17], PP1[17], PP2[17], PP3[17], PP4[17], PP5[17], PP6[17]);
  UB7_3C18 U14 (W0[20], W1[19], W2[18], PP0[18], PP1[18], PP2[18], PP3[18], PP4[18], PP5[18], PP6[18]);
  UB7_3C19 U15 (W0[21], W1[20], W2[19], PP0[19], PP1[19], PP2[19], PP3[19], PP4[19], PP5[19], PP6[19]);
  UB7_3C20 U16 (W0[22], W1[21], W2[20], PP0[20], PP1[20], PP2[20], PP3[20], PP4[20], PP5[20], PP6[20]);
  UB7_3C21 U17 (W0[23], W1[22], W2[21], PP0[21], PP1[21], PP2[21], PP3[21], PP4[21], PP5[21], PP6[21]);
  UB7_3C22 U18 (W0[24], W1[23], W2[22], PP0[22], PP1[22], PP2[22], PP3[22], PP4[22], PP5[22], PP6[22]);
  UB7_3C23 U19 (W0[25], W1[24], W2[23], PP0[23], PP1[23], PP2[23], PP3[23], PP4[23], PP5[23], PP6[23]);
  UB7_3C24 U20 (W0[26], W1[25], W2[24], PP0[24], PP1[24], PP2[24], PP3[24], PP4[24], PP5[24], PP6[24]);
  UB7_3C25 U21 (W0[27], W1[26], W2[25], PP0[25], PP1[25], PP2[25], PP3[25], PP4[25], PP5[25], PP6[25]);
  UB7_3C26 U22 (W0[28], W1[27], W2[26], PP0[26], PP1[26], PP2[26], PP3[26], PP4[26], PP5[26], PP6[26]);
  UB7_3C27 U23 (W0[29], W1[28], W2[27], PP0[27], PP1[27], PP2[27], PP3[27], PP4[27], PP5[27], PP6[27]);
  UB7_3C28 U24 (W0[30], W1[29], W2[28], PP0[28], PP1[28], PP2[28], PP3[28], PP4[28], PP5[28], PP6[28]);
  UB7_3C29 U25 (W0[31], W1[30], W2[29], PP0[29], PP1[29], PP2[29], PP3[29], PP4[29], PP5[29], PP6[29]);
  UB7_3C30 U26 (W0[32], W1[31], W2[30], PP0[30], PP1[30], PP2[30], PP3[30], PP4[30], PP5[30], PP6[30]);
  UB7_3C31 U27 (W0[33], W1[32], W2[31], PP0[31], PP1[31], PP2[31], PP3[31], PP4[31], PP5[31], PP6[31]);
  UB7_3C32 U28 (W0[34], W1[33], W2[32], PP0[32], PP1[32], PP2[32], PP3[32], PP4[32], PP5[32], PP6[32]);
  UB7_3C33 U29 (W0[35], W1[34], W2[33], PP0[33], PP1[33], PP2[33], PP3[33], PP4[33], PP5[33], PP6[33]);
  UB7_3C34 U30 (W0[36], W1[35], W2[34], PP0[34], PP1[34], PP2[34], PP3[34], PP4[34], PP5[34], PP6[34]);
  UB7_3C35 U31 (W0[37], W1[36], W2[35], PP0[35], PP1[35], PP2[35], PP3[35], PP4[35], PP5[35], PP6[35]);
  UB7_3C36 U32 (W0[38], W1[37], W2[36], PP0[36], PP1[36], PP2[36], PP3[36], PP4[36], PP5[36], PP6[36]);
  UB7_3C37 U33 (W0[39], W1[38], W2[37], PP0[37], PP1[37], PP2[37], PP3[37], PP4[37], PP5[37], PP6[37]);
  UB7_3C38 U34 (W0[40], W1[39], W2[38], PP0[38], PP1[38], PP2[38], PP3[38], PP4[38], PP5[38], PP6[38]);
  UB7_3C39 U35 (W0[41], W1[40], W2[39], PP0[39], PP1[39], PP2[39], PP3[39], PP4[39], PP5[39], PP6[39]);
  UB7_3C40 U36 (W0[42], W1[41], W2[40], PP0[40], PP1[40], PP2[40], PP3[40], PP4[40], PP5[40], PP6[40]);
  UB7_3C41 U37 (W0[43], W1[42], W2[41], PP0[41], PP1[41], PP2[41], PP3[41], PP4[41], PP5[41], PP6[41]);
  UB7_3C42 U38 (W0[44], W1[43], W2[42], PP0[42], PP1[42], PP2[42], PP3[42], PP4[42], PP5[42], PP6[42]);
  UB7_3C43 U39 (W0[45], W1[44], W2[43], PP0[43], PP1[43], PP2[43], PP3[43], PP4[43], PP5[43], PP6[43]);
  UB7_3C44 U40 (W0[46], W1[45], W2[44], PP0[44], PP1[44], PP2[44], PP3[44], PP4[44], PP5[44], PP6[44]);
  UB7_3C45 U41 (W0[47], W1[46], W2[45], PP0[45], PP1[45], PP2[45], PP3[45], PP4[45], PP5[45], PP6[45]);
  UB7_3C46 U42 (W0[48], W1[47], W2[46], PP0[46], PP1[46], PP2[46], PP3[46], PP4[46], PP5[46], PP6[46]);
  UB7_3C47 U43 (W0[49], W1[48], W2[47], PP0[47], PP1[47], PP2[47], PP3[47], PP4[47], PP5[47], PP6[47]);
  UB7_3C48 U44 (W0[50], W1[49], W2[48], PP0[48], PP1[48], PP2[48], PP3[48], PP4[48], PP5[48], PP6[48]);
  UB7_3C49 U45 (W0[51], W1[50], W2[49], PP0[49], PP1[49], PP2[49], PP3[49], PP4[49], PP5[49], PP6[49]);
  UB7_3C50 U46 (W0[52], W1[51], W2[50], PP0[50], PP1[50], PP2[50], PP3[50], PP4[50], PP5[50], PP6[50]);
  UB7_3C51 U47 (W0[53], W1[52], W2[51], PP0[51], PP1[51], PP2[51], PP3[51], PP4[51], PP5[51], PP6[51]);
  UB7_3C52 U48 (W0[54], W1[53], W2[52], PP0[52], PP1[52], PP2[52], PP3[52], PP4[52], PP5[52], PP6[52]);
  UB7_3C53 U49 (W0[55], W1[54], W2[53], PP0[53], PP1[53], PP2[53], PP3[53], PP4[53], PP5[53], PP6[53]);
  UB7_3C54 U50 (W0[56], W1[55], W2[54], PP0[54], PP1[54], PP2[54], PP3[54], PP4[54], PP5[54], PP6[54]);
  UB7_3C55 U51 (W0[57], W1[56], W2[55], PP0[55], PP1[55], PP2[55], PP3[55], PP4[55], PP5[55], PP6[55]);
  UB7_3C56 U52 (W0[58], W1[57], W2[56], PP0[56], PP1[56], PP2[56], PP3[56], PP4[56], PP5[56], PP6[56]);
  UB7_3C57 U53 (W0[59], W1[58], W2[57], PP0[57], PP1[57], PP2[57], PP3[57], PP4[57], PP5[57], PP6[57]);
  UB7_3C58 U54 (W0[60], W1[59], W2[58], PP0[58], PP1[58], PP2[58], PP3[58], PP4[58], PP5[58], PP6[58]);
  UB7_3C59 U55 (W0[61], W1[60], W2[59], PP0[59], PP1[59], PP2[59], PP3[59], PP4[59], PP5[59], PP6[59]);
  UB7_3C60 U56 (W0[62], W1[61], W2[60], PP0[60], PP1[60], PP2[60], PP3[60], PP4[60], PP5[60], PP6[60]);
  UB7_3C61 U57 (W0[63], W1[62], W2[61], PP0[61], PP1[61], PP2[61], PP3[61], PP4[61], PP5[61], PP6[61]);
  UB7_3C62 U58 (W0[64], W1[63], W2[62], PP0[62], PP1[62], PP2[62], PP3[62], PP4[62], PP5[62], PP6[62]);
  UB7_3C63 U59 (W0[65], W1[64], W2[63], PP0[63], PP1[63], PP2[63], PP3[63], PP4[63], PP5[63], PP6[63]);
  UB7_3C64 U60 (W0[66], W1[65], W2[64], PP0[64], PP1[64], PP2[64], PP3[64], PP4[64], PP5[64], PP6[64]);
  UB7_3C65 U61 (W0[67], W1[66], W2[65], PP0[65], PP1[65], PP2[65], PP3[65], PP4[65], PP5[65], PP6[65]);
  UB7_3C66 U62 (W0[68], W1[67], W2[66], PP0[66], PP1[66], PP2[66], PP3[66], PP4[66], PP5[66], PP6[66]);
  UB7_3C67 U63 (W0[69], W1[68], W2[67], PP0[67], PP1[67], PP2[67], PP3[67], PP4[67], PP5[67], PP6[67]);
  UB7_3C68 U64 (W0[70], W1[69], W2[68], PP0[68], PP1[68], PP2[68], PP3[68], PP4[68], PP5[68], PP6[68]);
  UB7_3C69 U65 (W0[71], W1[70], W2[69], PP0[69], PP1[69], PP2[69], PP3[69], PP4[69], PP5[69], PP6[69]);
  UB7_3C70 U66 (W0[72], W1[71], W2[70], PP0[70], PP1[70], PP2[70], PP3[70], PP4[70], PP5[70], PP6[70]);
  UB7_3C71 U67 (W0[73], W1[72], W2[71], PP0[71], PP1[71], PP2[71], PP3[71], PP4[71], PP5[71], PP6[71]);
  UB7_3C72 U68 (W0[74], W1[73], W2[72], PP0[72], PP1[72], PP2[72], PP3[72], PP4[72], PP5[72], PP6[72]);
  UB7_3C73 U69 (W0[75], W1[74], W2[73], PP0[73], PP1[73], PP2[73], PP3[73], PP4[73], PP5[73], PP6[73]);
  UB7_3C74 U70 (W0[76], W1[75], W2[74], PP0[74], PP1[74], PP2[74], PP3[74], PP4[74], PP5[74], PP6[74]);
  UB7_3C75 U71 (W0[77], W1[76], W2[75], PP0[75], PP1[75], PP2[75], PP3[75], PP4[75], PP5[75], PP6[75]);
  UB7_3C76 U72 (W0[78], W1[77], W2[76], PP0[76], PP1[76], PP2[76], PP3[76], PP4[76], PP5[76], PP6[76]);
  UB7_3C77 U73 (W0[79], W1[78], W2[77], PP0[77], PP1[77], PP2[77], PP3[77], PP4[77], PP5[77], PP6[77]);
  UB7_3C78 U74 (W0[80], W1[79], W2[78], PP0[78], PP1[78], PP2[78], PP3[78], PP4[78], PP5[78], PP6[78]);
  UB7_3C79 U75 (W0[81], W1[80], W2[79], PP0[79], PP1[79], PP2[79], PP3[79], PP4[79], PP5[79], PP6[79]);
  UB7_3C80 U76 (W0[82], W1[81], W2[80], PP0[80], PP1[80], PP2[80], PP3[80], PP4[80], PP5[80], PP6[80]);
  UB7_3C81 U77 (W0[83], W1[82], W2[81], PP0[81], PP1[81], PP2[81], PP3[81], PP4[81], PP5[81], PP6[81]);
  UB7_3C82 U78 (W0[84], W1[83], W2[82], PP0[82], PP1[82], PP2[82], PP3[82], PP4[82], PP5[82], PP6[82]);
  UB7_3C83 U79 (W0[85], W1[84], W2[83], PP0[83], PP1[83], PP2[83], PP3[83], PP4[83], PP5[83], PP6[83]);
  UB7_3C84 U80 (W0[86], W1[85], W2[84], PP0[84], PP1[84], PP2[84], PP3[84], PP4[84], PP5[84], PP6[84]);
  UB7_3C85 U81 (W0[87], W1[86], W2[85], PP0[85], PP1[85], PP2[85], PP3[85], PP4[85], PP5[85], PP6[85]);
  UB7_3C86 U82 (W0[88], W1[87], W2[86], PP0[86], PP1[86], PP2[86], PP3[86], PP4[86], PP5[86], PP6[86]);
  UB7_3C87 U83 (W0[89], W1[88], W2[87], PP0[87], PP1[87], PP2[87], PP3[87], PP4[87], PP5[87], PP6[87]);
  UB7_3C88 U84 (W0[90], W1[89], W2[88], PP0[88], PP1[88], PP2[88], PP3[88], PP4[88], PP5[88], PP6[88]);
  UB7_3C89 U85 (W0[91], W1[90], W2[89], PP0[89], PP1[89], PP2[89], PP3[89], PP4[89], PP5[89], PP6[89]);
  UB7_3C90 U86 (W0[92], W1[91], W2[90], PP0[90], PP1[90], PP2[90], PP3[90], PP4[90], PP5[90], PP6[90]);
  UB7_3C91 U87 (W0[93], W1[92], W2[91], PP0[91], PP1[91], PP2[91], PP3[91], PP4[91], PP5[91], PP6[91]);
  UB7_3C92 U88 (W0[94], W1[93], W2[92], PP0[92], PP1[92], PP2[92], PP3[92], PP4[92], PP5[92], PP6[92]);
  UB7_3C93 U89 (W0[95], W1[94], W2[93], PP0[93], PP1[93], PP2[93], PP3[93], PP4[93], PP5[93], PP6[93]);
  UB7_3C94 U90 (W0[96], W1[95], W2[94], PP0[94], PP1[94], PP2[94], PP3[94], PP4[94], PP5[94], PP6[94]);
  UB7_3C95 U91 (W0[97], W1[96], W2[95], PP0[95], PP1[95], PP2[95], PP3[95], PP4[95], PP5[95], PP6[95]);
  UB7_3C96 U92 (W0[98], W1[97], W2[96], PP0[96], PP1[96], PP2[96], PP3[96], PP4[96], PP5[96], PP6[96]);
  UB7_3C97 U93 (W0[99], W1[98], W2[97], PP0[97], PP1[97], PP2[97], PP3[97], PP4[97], PP5[97], PP6[97]);
  UB7_3C98 U94 (W0[100], W1[99], W2[98], PP0[98], PP1[98], PP2[98], PP3[98], PP4[98], PP5[98], PP6[98]);
  UB7_3C99 U95 (W0[101], W1[100], W2[99], PP0[99], PP1[99], PP2[99], PP3[99], PP4[99], PP5[99], PP6[99]);
  UB7_3C100 U96 (W0[102], W1[101], W2[100], PP0[100], PP1[100], PP2[100], PP3[100], PP4[100], PP5[100], PP6[100]);
  UB7_3C101 U97 (W0[103], W1[102], W2[101], PP0[101], PP1[101], PP2[101], PP3[101], PP4[101], PP5[101], PP6[101]);
  UB7_3C102 U98 (W0[104], W1[103], W2[102], PP0[102], PP1[102], PP2[102], PP3[102], PP4[102], PP5[102], PP6[102]);
  UB7_3C103 U99 (W0[105], W1[104], W2[103], PP0[103], PP1[103], PP2[103], PP3[103], PP4[103], PP5[103], PP6[103]);
  UB7_3C104 U100 (W0[106], W1[105], W2[104], PP0[104], PP1[104], PP2[104], PP3[104], PP4[104], PP5[104], PP6[104]);
  UB7_3C105 U101 (W0[107], W1[106], W2[105], PP0[105], PP1[105], PP2[105], PP3[105], PP4[105], PP5[105], PP6[105]);
  UB7_3C106 U102 (W0[108], W1[107], W2[106], PP0[106], PP1[106], PP2[106], PP3[106], PP4[106], PP5[106], PP6[106]);
  UB7_3C107 U103 (W0[109], W1[108], W2[107], PP0[107], PP1[107], PP2[107], PP3[107], PP4[107], PP5[107], PP6[107]);
  UB7_3C108 U104 (W0[110], W1[109], W2[108], PP0[108], PP1[108], PP2[108], PP3[108], PP4[108], PP5[108], PP6[108]);
  UB7_3C109 U105 (W0[111], W1[110], W2[109], PP0[109], PP1[109], PP2[109], PP3[109], PP4[109], PP5[109], PP6[109]);
  UB7_3C110 U106 (W0[112], W1[111], W2[110], PP0[110], PP1[110], PP2[110], PP3[110], PP4[110], PP5[110], PP6[110]);
  UB7_3C111 U107 (W0[113], W1[112], W2[111], PP0[111], PP1[111], PP2[111], PP3[111], PP4[111], PP5[111], PP6[111]);
  UB7_3C112 U108 (W0[114], W1[113], W2[112], PP0[112], PP1[112], PP2[112], PP3[112], PP4[112], PP5[112], PP6[112]);
  UB7_3C113 U109 (W0[115], W1[114], W2[113], PP0[113], PP1[113], PP2[113], PP3[113], PP4[113], PP5[113], PP6[113]);
  UB7_3C114 U110 (W0[116], W1[115], W2[114], PP0[114], PP1[114], PP2[114], PP3[114], PP4[114], PP5[114], PP6[114]);
  UB7_3C115 U111 (W0[117], W1[116], W2[115], PP0[115], PP1[115], PP2[115], PP3[115], PP4[115], PP5[115], PP6[115]);
  UB7_3C116 U112 (W0[118], W1[117], W2[116], PP0[116], PP1[116], PP2[116], PP3[116], PP4[116], PP5[116], PP6[116]);
  UB6_3C117 U113 (W0[119], W1[118], W2[117], PP0[117], PP1[117], PP2[117], PP3[117], PP4[117], PP5[117]);
  UB5_3C118 U114 (W0[120], W1[119], W2[118], PP0[118], PP1[118], PP2[118], PP3[118], PP4[118]);
  UB5_3C119 U115 (W0[121], W1[120], W2[119], PP0[119], PP1[119], PP2[119], PP3[119], PP4[119]);
  UB4_3C120 U116 (W0[122], W1[121], W2[120], PP0[120], PP1[120], PP2[120], PP3[120]);
  UB4_3C121 U117 (W0[123], W1[122], W2[121], PP0[121], PP1[121], PP2[121], PP3[121]);
  UBFA_122 U118 (W1[123], W2[122], PP0[122], PP1[122], PP2[122]);
  UBFA_123 U119 (W2[124], W2[123], PP0[123], PP1[123], PP2[123]);
  UBCON_3_0 U120 (W0[3:0], PP0[3:0]);
  UB1DCON_4 U121 (W0[4], PP2[4]);
  UB1DCON_5 U122 (W0[5], PP3[5]);
  UBCON_7_6 U123 (W0[7:6], PP4[7:6]);
  UBCON_126_124 U124 (W0[126:124], PP0[126:124]);
  UBCON_3_0 U125 (W1[3:0], PP1[3:0]);
  UB1DCON_4 U126 (W1[4], PP3[4]);
  UBCON_125_124 U127 (W1[125:124], PP1[125:124]);
  UBCON_3_2 U128 (W2[3:2], PP2[3:2]);
  D7_3CTR_126_0_125002 U129 (S1, S2, W0, W1, W2);
endmodule

module D7_3CTR_126_0_125002 (S1, S2, PP0, PP1, PP2);
  output [126:0] S1;
  output [126:0] S2;
  input [126:0] PP0;
  input [125:0] PP1;
  input [124:2] PP2;
  wire [126:0] W0;
  wire [126:0] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W0[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U10 (W0[13], W1[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U11 (W0[14], W1[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U12 (W0[15], W1[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U13 (W0[16], W1[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U14 (W0[17], W1[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U15 (W0[18], W1[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U16 (W0[19], W1[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U17 (W0[20], W1[19], PP0[19], PP1[19], PP2[19]);
  UBFA_20 U18 (W0[21], W1[20], PP0[20], PP1[20], PP2[20]);
  UBFA_21 U19 (W0[22], W1[21], PP0[21], PP1[21], PP2[21]);
  UBFA_22 U20 (W0[23], W1[22], PP0[22], PP1[22], PP2[22]);
  UBFA_23 U21 (W0[24], W1[23], PP0[23], PP1[23], PP2[23]);
  UBFA_24 U22 (W0[25], W1[24], PP0[24], PP1[24], PP2[24]);
  UBFA_25 U23 (W0[26], W1[25], PP0[25], PP1[25], PP2[25]);
  UBFA_26 U24 (W0[27], W1[26], PP0[26], PP1[26], PP2[26]);
  UBFA_27 U25 (W0[28], W1[27], PP0[27], PP1[27], PP2[27]);
  UBFA_28 U26 (W0[29], W1[28], PP0[28], PP1[28], PP2[28]);
  UBFA_29 U27 (W0[30], W1[29], PP0[29], PP1[29], PP2[29]);
  UBFA_30 U28 (W0[31], W1[30], PP0[30], PP1[30], PP2[30]);
  UBFA_31 U29 (W0[32], W1[31], PP0[31], PP1[31], PP2[31]);
  UBFA_32 U30 (W0[33], W1[32], PP0[32], PP1[32], PP2[32]);
  UBFA_33 U31 (W0[34], W1[33], PP0[33], PP1[33], PP2[33]);
  UBFA_34 U32 (W0[35], W1[34], PP0[34], PP1[34], PP2[34]);
  UBFA_35 U33 (W0[36], W1[35], PP0[35], PP1[35], PP2[35]);
  UBFA_36 U34 (W0[37], W1[36], PP0[36], PP1[36], PP2[36]);
  UBFA_37 U35 (W0[38], W1[37], PP0[37], PP1[37], PP2[37]);
  UBFA_38 U36 (W0[39], W1[38], PP0[38], PP1[38], PP2[38]);
  UBFA_39 U37 (W0[40], W1[39], PP0[39], PP1[39], PP2[39]);
  UBFA_40 U38 (W0[41], W1[40], PP0[40], PP1[40], PP2[40]);
  UBFA_41 U39 (W0[42], W1[41], PP0[41], PP1[41], PP2[41]);
  UBFA_42 U40 (W0[43], W1[42], PP0[42], PP1[42], PP2[42]);
  UBFA_43 U41 (W0[44], W1[43], PP0[43], PP1[43], PP2[43]);
  UBFA_44 U42 (W0[45], W1[44], PP0[44], PP1[44], PP2[44]);
  UBFA_45 U43 (W0[46], W1[45], PP0[45], PP1[45], PP2[45]);
  UBFA_46 U44 (W0[47], W1[46], PP0[46], PP1[46], PP2[46]);
  UBFA_47 U45 (W0[48], W1[47], PP0[47], PP1[47], PP2[47]);
  UBFA_48 U46 (W0[49], W1[48], PP0[48], PP1[48], PP2[48]);
  UBFA_49 U47 (W0[50], W1[49], PP0[49], PP1[49], PP2[49]);
  UBFA_50 U48 (W0[51], W1[50], PP0[50], PP1[50], PP2[50]);
  UBFA_51 U49 (W0[52], W1[51], PP0[51], PP1[51], PP2[51]);
  UBFA_52 U50 (W0[53], W1[52], PP0[52], PP1[52], PP2[52]);
  UBFA_53 U51 (W0[54], W1[53], PP0[53], PP1[53], PP2[53]);
  UBFA_54 U52 (W0[55], W1[54], PP0[54], PP1[54], PP2[54]);
  UBFA_55 U53 (W0[56], W1[55], PP0[55], PP1[55], PP2[55]);
  UBFA_56 U54 (W0[57], W1[56], PP0[56], PP1[56], PP2[56]);
  UBFA_57 U55 (W0[58], W1[57], PP0[57], PP1[57], PP2[57]);
  UBFA_58 U56 (W0[59], W1[58], PP0[58], PP1[58], PP2[58]);
  UBFA_59 U57 (W0[60], W1[59], PP0[59], PP1[59], PP2[59]);
  UBFA_60 U58 (W0[61], W1[60], PP0[60], PP1[60], PP2[60]);
  UBFA_61 U59 (W0[62], W1[61], PP0[61], PP1[61], PP2[61]);
  UBFA_62 U60 (W0[63], W1[62], PP0[62], PP1[62], PP2[62]);
  UBFA_63 U61 (W0[64], W1[63], PP0[63], PP1[63], PP2[63]);
  UBFA_64 U62 (W0[65], W1[64], PP0[64], PP1[64], PP2[64]);
  UBFA_65 U63 (W0[66], W1[65], PP0[65], PP1[65], PP2[65]);
  UBFA_66 U64 (W0[67], W1[66], PP0[66], PP1[66], PP2[66]);
  UBFA_67 U65 (W0[68], W1[67], PP0[67], PP1[67], PP2[67]);
  UBFA_68 U66 (W0[69], W1[68], PP0[68], PP1[68], PP2[68]);
  UBFA_69 U67 (W0[70], W1[69], PP0[69], PP1[69], PP2[69]);
  UBFA_70 U68 (W0[71], W1[70], PP0[70], PP1[70], PP2[70]);
  UBFA_71 U69 (W0[72], W1[71], PP0[71], PP1[71], PP2[71]);
  UBFA_72 U70 (W0[73], W1[72], PP0[72], PP1[72], PP2[72]);
  UBFA_73 U71 (W0[74], W1[73], PP0[73], PP1[73], PP2[73]);
  UBFA_74 U72 (W0[75], W1[74], PP0[74], PP1[74], PP2[74]);
  UBFA_75 U73 (W0[76], W1[75], PP0[75], PP1[75], PP2[75]);
  UBFA_76 U74 (W0[77], W1[76], PP0[76], PP1[76], PP2[76]);
  UBFA_77 U75 (W0[78], W1[77], PP0[77], PP1[77], PP2[77]);
  UBFA_78 U76 (W0[79], W1[78], PP0[78], PP1[78], PP2[78]);
  UBFA_79 U77 (W0[80], W1[79], PP0[79], PP1[79], PP2[79]);
  UBFA_80 U78 (W0[81], W1[80], PP0[80], PP1[80], PP2[80]);
  UBFA_81 U79 (W0[82], W1[81], PP0[81], PP1[81], PP2[81]);
  UBFA_82 U80 (W0[83], W1[82], PP0[82], PP1[82], PP2[82]);
  UBFA_83 U81 (W0[84], W1[83], PP0[83], PP1[83], PP2[83]);
  UBFA_84 U82 (W0[85], W1[84], PP0[84], PP1[84], PP2[84]);
  UBFA_85 U83 (W0[86], W1[85], PP0[85], PP1[85], PP2[85]);
  UBFA_86 U84 (W0[87], W1[86], PP0[86], PP1[86], PP2[86]);
  UBFA_87 U85 (W0[88], W1[87], PP0[87], PP1[87], PP2[87]);
  UBFA_88 U86 (W0[89], W1[88], PP0[88], PP1[88], PP2[88]);
  UBFA_89 U87 (W0[90], W1[89], PP0[89], PP1[89], PP2[89]);
  UBFA_90 U88 (W0[91], W1[90], PP0[90], PP1[90], PP2[90]);
  UBFA_91 U89 (W0[92], W1[91], PP0[91], PP1[91], PP2[91]);
  UBFA_92 U90 (W0[93], W1[92], PP0[92], PP1[92], PP2[92]);
  UBFA_93 U91 (W0[94], W1[93], PP0[93], PP1[93], PP2[93]);
  UBFA_94 U92 (W0[95], W1[94], PP0[94], PP1[94], PP2[94]);
  UBFA_95 U93 (W0[96], W1[95], PP0[95], PP1[95], PP2[95]);
  UBFA_96 U94 (W0[97], W1[96], PP0[96], PP1[96], PP2[96]);
  UBFA_97 U95 (W0[98], W1[97], PP0[97], PP1[97], PP2[97]);
  UBFA_98 U96 (W0[99], W1[98], PP0[98], PP1[98], PP2[98]);
  UBFA_99 U97 (W0[100], W1[99], PP0[99], PP1[99], PP2[99]);
  UBFA_100 U98 (W0[101], W1[100], PP0[100], PP1[100], PP2[100]);
  UBFA_101 U99 (W0[102], W1[101], PP0[101], PP1[101], PP2[101]);
  UBFA_102 U100 (W0[103], W1[102], PP0[102], PP1[102], PP2[102]);
  UBFA_103 U101 (W0[104], W1[103], PP0[103], PP1[103], PP2[103]);
  UBFA_104 U102 (W0[105], W1[104], PP0[104], PP1[104], PP2[104]);
  UBFA_105 U103 (W0[106], W1[105], PP0[105], PP1[105], PP2[105]);
  UBFA_106 U104 (W0[107], W1[106], PP0[106], PP1[106], PP2[106]);
  UBFA_107 U105 (W0[108], W1[107], PP0[107], PP1[107], PP2[107]);
  UBFA_108 U106 (W0[109], W1[108], PP0[108], PP1[108], PP2[108]);
  UBFA_109 U107 (W0[110], W1[109], PP0[109], PP1[109], PP2[109]);
  UBFA_110 U108 (W0[111], W1[110], PP0[110], PP1[110], PP2[110]);
  UBFA_111 U109 (W0[112], W1[111], PP0[111], PP1[111], PP2[111]);
  UBFA_112 U110 (W0[113], W1[112], PP0[112], PP1[112], PP2[112]);
  UBFA_113 U111 (W0[114], W1[113], PP0[113], PP1[113], PP2[113]);
  UBFA_114 U112 (W0[115], W1[114], PP0[114], PP1[114], PP2[114]);
  UBFA_115 U113 (W0[116], W1[115], PP0[115], PP1[115], PP2[115]);
  UBFA_116 U114 (W0[117], W1[116], PP0[116], PP1[116], PP2[116]);
  UBFA_117 U115 (W0[118], W1[117], PP0[117], PP1[117], PP2[117]);
  UBFA_118 U116 (W0[119], W1[118], PP0[118], PP1[118], PP2[118]);
  UBFA_119 U117 (W0[120], W1[119], PP0[119], PP1[119], PP2[119]);
  UBFA_120 U118 (W0[121], W1[120], PP0[120], PP1[120], PP2[120]);
  UBFA_121 U119 (W0[122], W1[121], PP0[121], PP1[121], PP2[121]);
  UBFA_122 U120 (W0[123], W1[122], PP0[122], PP1[122], PP2[122]);
  UBFA_123 U121 (W0[124], W1[123], PP0[123], PP1[123], PP2[123]);
  UBFA_124 U122 (W0[125], W1[124], PP0[124], PP1[124], PP2[124]);
  UBHA_125 U123 (W1[126], W1[125], PP0[125], PP1[125]);
  UBCON_1_0 U124 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U125 (W0[2], PP2[2]);
  UB1DCON_126 U126 (W0[126], PP0[126]);
  UBCON_1_0 U127 (W1[1:0], PP1[1:0]);
  D7_3CTR_126_0_126000 U128 (S1, S2, W0, W1);
endmodule

module D7_3CTR_126_0_126000 (S1, S2, PP0, PP1);
  output [126:0] S1;
  output [126:0] S2;
  input [126:0] PP0;
  input [126:0] PP1;
  UBCON_126_0 U0 (S1, PP0);
  UBCON_126_0 U1 (S2, PP1);
endmodule

module D7_3CTR_65_0_67_0000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, PP32);
  output [126:0] S1;
  output [126:0] S2;
  input [65:0] PP0;
  input [67:0] PP1;
  input [85:18] PP10;
  input [87:20] PP11;
  input [89:22] PP12;
  input [91:24] PP13;
  input [93:26] PP14;
  input [95:28] PP15;
  input [97:30] PP16;
  input [99:32] PP17;
  input [101:34] PP18;
  input [103:36] PP19;
  input [69:2] PP2;
  input [105:38] PP20;
  input [107:40] PP21;
  input [109:42] PP22;
  input [111:44] PP23;
  input [113:46] PP24;
  input [115:48] PP25;
  input [117:50] PP26;
  input [119:52] PP27;
  input [121:54] PP28;
  input [123:56] PP29;
  input [71:4] PP3;
  input [125:58] PP30;
  input [126:60] PP31;
  input [64:62] PP32;
  input [73:6] PP4;
  input [75:8] PP5;
  input [77:10] PP6;
  input [79:12] PP7;
  input [81:14] PP8;
  input [83:16] PP9;
  wire [126:0] W0;
  wire [125:0] W1;
  wire [107:18] W10;
  wire [105:20] W11;
  wire [103:22] W12;
  wire [101:24] W13;
  wire [100:26] W14;
  wire [123:2] W2;
  wire [121:4] W3;
  wire [119:6] W4;
  wire [117:8] W5;
  wire [115:10] W6;
  wire [113:12] W7;
  wire [111:14] W8;
  wire [109:16] W9;
  UBHA_28 U0 (W13[29], W14[28], PP0[28], PP1[28]);
  UBFA_29 U1 (W13[30], W14[29], PP0[29], PP1[29], PP2[29]);
  UB4_3C30 U2 (W12[32], W13[31], W14[30], PP0[30], PP1[30], PP2[30], PP3[30]);
  UB4_3C31 U3 (W12[33], W13[32], W14[31], PP0[31], PP1[31], PP2[31], PP3[31]);
  UB6_3C32 U4 (W12[34], W13[33], W14[32], PP0[32], PP1[32], PP2[32], PP3[32], PP4[32], PP5[32]);
  UB6_3C33 U5 (W12[35], W13[34], W14[33], PP0[33], PP1[33], PP2[33], PP3[33], PP4[33], PP5[33]);
  UB7_3C34 U6 (W11[36], W13[35], W14[34], PP0[34], PP1[34], PP2[34], PP3[34], PP4[34], PP5[34], PP6[34]);
  UB7_3C35 U7 (W10[37], W12[36], W14[35], PP0[35], PP1[35], PP2[35], PP3[35], PP4[35], PP5[35], PP6[35]);
  UB7_3C36 U8 (W10[38], W11[37], W13[36], PP0[36], PP1[36], PP2[36], PP3[36], PP4[36], PP5[36], PP6[36]);
  UBHA_36 U9 (W12[37], W14[36], PP7[36], PP8[36]);
  UB7_3C37 U10 (W10[39], W11[38], W13[37], PP0[37], PP1[37], PP2[37], PP3[37], PP4[37], PP5[37], PP6[37]);
  UBFA_37 U11 (W12[38], W14[37], PP7[37], PP8[37], PP9[37]);
  UB7_3C38 U12 (W9[40], W11[39], W13[38], PP0[38], PP1[38], PP2[38], PP3[38], PP4[38], PP5[38], PP6[38]);
  UB4_3C38 U13 (W10[40], W12[39], W14[38], PP7[38], PP8[38], PP9[38], PP10[38]);
  UB7_3C39 U14 (W9[41], W11[40], W13[39], PP0[39], PP1[39], PP2[39], PP3[39], PP4[39], PP5[39], PP6[39]);
  UB4_3C39 U15 (W10[41], W12[40], W14[39], PP7[39], PP8[39], PP9[39], PP10[39]);
  UB7_3C40 U16 (W9[42], W11[41], W13[40], PP0[40], PP1[40], PP2[40], PP3[40], PP4[40], PP5[40], PP6[40]);
  UB6_3C40 U17 (W10[42], W12[41], W14[40], PP7[40], PP8[40], PP9[40], PP10[40], PP11[40], PP12[40]);
  UB7_3C41 U18 (W9[43], W11[42], W13[41], PP0[41], PP1[41], PP2[41], PP3[41], PP4[41], PP5[41], PP6[41]);
  UB6_3C41 U19 (W10[43], W12[42], W14[41], PP7[41], PP8[41], PP9[41], PP10[41], PP11[41], PP12[41]);
  UB7_3C42 U20 (W8[44], W11[43], W13[42], PP0[42], PP1[42], PP2[42], PP3[42], PP4[42], PP5[42], PP6[42]);
  UB7_3C42 U21 (W9[44], W12[43], W14[42], PP7[42], PP8[42], PP9[42], PP10[42], PP11[42], PP12[42], PP13[42]);
  UB7_3C43 U22 (W7[45], W10[44], W13[43], PP0[43], PP1[43], PP2[43], PP3[43], PP4[43], PP5[43], PP6[43]);
  UB7_3C43 U23 (W8[45], W11[44], W14[43], PP7[43], PP8[43], PP9[43], PP10[43], PP11[43], PP12[43], PP13[43]);
  UB7_3C44 U24 (W7[46], W9[45], W12[44], PP0[44], PP1[44], PP2[44], PP3[44], PP4[44], PP5[44], PP6[44]);
  UB7_3C44 U25 (W8[46], W10[45], W13[44], PP7[44], PP8[44], PP9[44], PP10[44], PP11[44], PP12[44], PP13[44]);
  UBHA_44 U26 (W11[45], W14[44], PP14[44], PP15[44]);
  UB7_3C45 U27 (W7[47], W9[46], W12[45], PP0[45], PP1[45], PP2[45], PP3[45], PP4[45], PP5[45], PP6[45]);
  UB7_3C45 U28 (W8[47], W10[46], W13[45], PP7[45], PP8[45], PP9[45], PP10[45], PP11[45], PP12[45], PP13[45]);
  UBFA_45 U29 (W11[46], W14[45], PP14[45], PP15[45], PP16[45]);
  UB7_3C46 U30 (W6[48], W9[47], W12[46], PP0[46], PP1[46], PP2[46], PP3[46], PP4[46], PP5[46], PP6[46]);
  UB7_3C46 U31 (W7[48], W10[47], W13[46], PP7[46], PP8[46], PP9[46], PP10[46], PP11[46], PP12[46], PP13[46]);
  UB4_3C46 U32 (W8[48], W11[47], W14[46], PP14[46], PP15[46], PP16[46], PP17[46]);
  UB7_3C47 U33 (W6[49], W9[48], W12[47], PP0[47], PP1[47], PP2[47], PP3[47], PP4[47], PP5[47], PP6[47]);
  UB7_3C47 U34 (W7[49], W10[48], W13[47], PP7[47], PP8[47], PP9[47], PP10[47], PP11[47], PP12[47], PP13[47]);
  UB4_3C47 U35 (W8[49], W11[48], W14[47], PP14[47], PP15[47], PP16[47], PP17[47]);
  UB7_3C48 U36 (W6[50], W9[49], W12[48], PP0[48], PP1[48], PP2[48], PP3[48], PP4[48], PP5[48], PP6[48]);
  UB7_3C48 U37 (W7[50], W10[49], W13[48], PP7[48], PP8[48], PP9[48], PP10[48], PP11[48], PP12[48], PP13[48]);
  UB6_3C48 U38 (W8[50], W11[49], W14[48], PP14[48], PP15[48], PP16[48], PP17[48], PP18[48], PP19[48]);
  UB7_3C49 U39 (W6[51], W9[50], W12[49], PP0[49], PP1[49], PP2[49], PP3[49], PP4[49], PP5[49], PP6[49]);
  UB7_3C49 U40 (W7[51], W10[50], W13[49], PP7[49], PP8[49], PP9[49], PP10[49], PP11[49], PP12[49], PP13[49]);
  UB6_3C49 U41 (W8[51], W11[50], W14[49], PP14[49], PP15[49], PP16[49], PP17[49], PP18[49], PP19[49]);
  UB7_3C50 U42 (W5[52], W9[51], W12[50], PP0[50], PP1[50], PP2[50], PP3[50], PP4[50], PP5[50], PP6[50]);
  UB7_3C50 U43 (W6[52], W10[51], W13[50], PP7[50], PP8[50], PP9[50], PP10[50], PP11[50], PP12[50], PP13[50]);
  UB7_3C50 U44 (W7[52], W11[51], W14[50], PP14[50], PP15[50], PP16[50], PP17[50], PP18[50], PP19[50], PP20[50]);
  UB7_3C51 U45 (W4[53], W8[52], W12[51], PP0[51], PP1[51], PP2[51], PP3[51], PP4[51], PP5[51], PP6[51]);
  UB7_3C51 U46 (W5[53], W9[52], W13[51], PP7[51], PP8[51], PP9[51], PP10[51], PP11[51], PP12[51], PP13[51]);
  UB7_3C51 U47 (W6[53], W10[52], W14[51], PP14[51], PP15[51], PP16[51], PP17[51], PP18[51], PP19[51], PP20[51]);
  UB7_3C52 U48 (W4[54], W7[53], W11[52], PP0[52], PP1[52], PP2[52], PP3[52], PP4[52], PP5[52], PP6[52]);
  UB7_3C52 U49 (W5[54], W8[53], W12[52], PP7[52], PP8[52], PP9[52], PP10[52], PP11[52], PP12[52], PP13[52]);
  UB7_3C52 U50 (W6[54], W9[53], W13[52], PP14[52], PP15[52], PP16[52], PP17[52], PP18[52], PP19[52], PP20[52]);
  UBHA_52 U51 (W10[53], W14[52], PP21[52], PP22[52]);
  UB7_3C53 U52 (W4[55], W7[54], W11[53], PP0[53], PP1[53], PP2[53], PP3[53], PP4[53], PP5[53], PP6[53]);
  UB7_3C53 U53 (W5[55], W8[54], W12[53], PP7[53], PP8[53], PP9[53], PP10[53], PP11[53], PP12[53], PP13[53]);
  UB7_3C53 U54 (W6[55], W9[54], W13[53], PP14[53], PP15[53], PP16[53], PP17[53], PP18[53], PP19[53], PP20[53]);
  UBFA_53 U55 (W10[54], W14[53], PP21[53], PP22[53], PP23[53]);
  UB7_3C54 U56 (W3[56], W7[55], W11[54], PP0[54], PP1[54], PP2[54], PP3[54], PP4[54], PP5[54], PP6[54]);
  UB7_3C54 U57 (W4[56], W8[55], W12[54], PP7[54], PP8[54], PP9[54], PP10[54], PP11[54], PP12[54], PP13[54]);
  UB7_3C54 U58 (W5[56], W9[55], W13[54], PP14[54], PP15[54], PP16[54], PP17[54], PP18[54], PP19[54], PP20[54]);
  UB4_3C54 U59 (W6[56], W10[55], W14[54], PP21[54], PP22[54], PP23[54], PP24[54]);
  UB7_3C55 U60 (W3[57], W7[56], W11[55], PP0[55], PP1[55], PP2[55], PP3[55], PP4[55], PP5[55], PP6[55]);
  UB7_3C55 U61 (W4[57], W8[56], W12[55], PP7[55], PP8[55], PP9[55], PP10[55], PP11[55], PP12[55], PP13[55]);
  UB7_3C55 U62 (W5[57], W9[56], W13[55], PP14[55], PP15[55], PP16[55], PP17[55], PP18[55], PP19[55], PP20[55]);
  UB4_3C55 U63 (W6[57], W10[56], W14[55], PP21[55], PP22[55], PP23[55], PP24[55]);
  UB7_3C56 U64 (W3[58], W7[57], W11[56], PP0[56], PP1[56], PP2[56], PP3[56], PP4[56], PP5[56], PP6[56]);
  UB7_3C56 U65 (W4[58], W8[57], W12[56], PP7[56], PP8[56], PP9[56], PP10[56], PP11[56], PP12[56], PP13[56]);
  UB7_3C56 U66 (W5[58], W9[57], W13[56], PP14[56], PP15[56], PP16[56], PP17[56], PP18[56], PP19[56], PP20[56]);
  UB6_3C56 U67 (W6[58], W10[57], W14[56], PP21[56], PP22[56], PP23[56], PP24[56], PP25[56], PP26[56]);
  UB7_3C57 U68 (W3[59], W7[58], W11[57], PP0[57], PP1[57], PP2[57], PP3[57], PP4[57], PP5[57], PP6[57]);
  UB7_3C57 U69 (W4[59], W8[58], W12[57], PP7[57], PP8[57], PP9[57], PP10[57], PP11[57], PP12[57], PP13[57]);
  UB7_3C57 U70 (W5[59], W9[58], W13[57], PP14[57], PP15[57], PP16[57], PP17[57], PP18[57], PP19[57], PP20[57]);
  UB6_3C57 U71 (W6[59], W10[58], W14[57], PP21[57], PP22[57], PP23[57], PP24[57], PP25[57], PP26[57]);
  UB7_3C58 U72 (W2[60], W7[59], W11[58], PP0[58], PP1[58], PP2[58], PP3[58], PP4[58], PP5[58], PP6[58]);
  UB7_3C58 U73 (W3[60], W8[59], W12[58], PP7[58], PP8[58], PP9[58], PP10[58], PP11[58], PP12[58], PP13[58]);
  UB7_3C58 U74 (W4[60], W9[59], W13[58], PP14[58], PP15[58], PP16[58], PP17[58], PP18[58], PP19[58], PP20[58]);
  UB7_3C58 U75 (W5[60], W10[59], W14[58], PP21[58], PP22[58], PP23[58], PP24[58], PP25[58], PP26[58], PP27[58]);
  UB7_3C59 U76 (W1[61], W6[60], W11[59], PP0[59], PP1[59], PP2[59], PP3[59], PP4[59], PP5[59], PP6[59]);
  UB7_3C59 U77 (W2[61], W7[60], W12[59], PP7[59], PP8[59], PP9[59], PP10[59], PP11[59], PP12[59], PP13[59]);
  UB7_3C59 U78 (W3[61], W8[60], W13[59], PP14[59], PP15[59], PP16[59], PP17[59], PP18[59], PP19[59], PP20[59]);
  UB7_3C59 U79 (W4[61], W9[60], W14[59], PP21[59], PP22[59], PP23[59], PP24[59], PP25[59], PP26[59], PP27[59]);
  UB7_3C60 U80 (W1[62], W5[61], W10[60], PP0[60], PP1[60], PP2[60], PP3[60], PP4[60], PP5[60], PP6[60]);
  UB7_3C60 U81 (W2[62], W6[61], W11[60], PP7[60], PP8[60], PP9[60], PP10[60], PP11[60], PP12[60], PP13[60]);
  UB7_3C60 U82 (W3[62], W7[61], W12[60], PP14[60], PP15[60], PP16[60], PP17[60], PP18[60], PP19[60], PP20[60]);
  UB7_3C60 U83 (W4[62], W8[61], W13[60], PP21[60], PP22[60], PP23[60], PP24[60], PP25[60], PP26[60], PP27[60]);
  UBHA_60 U84 (W9[61], W14[60], PP28[60], PP29[60]);
  UB7_3C61 U85 (W1[63], W5[62], W10[61], PP0[61], PP1[61], PP2[61], PP3[61], PP4[61], PP5[61], PP6[61]);
  UB7_3C61 U86 (W2[63], W6[62], W11[61], PP7[61], PP8[61], PP9[61], PP10[61], PP11[61], PP12[61], PP13[61]);
  UB7_3C61 U87 (W3[63], W7[62], W12[61], PP14[61], PP15[61], PP16[61], PP17[61], PP18[61], PP19[61], PP20[61]);
  UB7_3C61 U88 (W4[63], W8[62], W13[61], PP21[61], PP22[61], PP23[61], PP24[61], PP25[61], PP26[61], PP27[61]);
  UBFA_61 U89 (W9[62], W14[61], PP28[61], PP29[61], PP30[61]);
  UB7_3C62 U90 (W0[64], W5[63], W10[62], PP0[62], PP1[62], PP2[62], PP3[62], PP4[62], PP5[62], PP6[62]);
  UB7_3C62 U91 (W1[64], W6[63], W11[62], PP7[62], PP8[62], PP9[62], PP10[62], PP11[62], PP12[62], PP13[62]);
  UB7_3C62 U92 (W2[64], W7[63], W12[62], PP14[62], PP15[62], PP16[62], PP17[62], PP18[62], PP19[62], PP20[62]);
  UB7_3C62 U93 (W3[64], W8[63], W13[62], PP21[62], PP22[62], PP23[62], PP24[62], PP25[62], PP26[62], PP27[62]);
  UB4_3C62 U94 (W4[64], W9[63], W14[62], PP28[62], PP29[62], PP30[62], PP31[62]);
  UB7_3C63 U95 (W0[65], W5[64], W10[63], PP0[63], PP1[63], PP2[63], PP3[63], PP4[63], PP5[63], PP6[63]);
  UB7_3C63 U96 (W1[65], W6[64], W11[63], PP7[63], PP8[63], PP9[63], PP10[63], PP11[63], PP12[63], PP13[63]);
  UB7_3C63 U97 (W2[65], W7[64], W12[63], PP14[63], PP15[63], PP16[63], PP17[63], PP18[63], PP19[63], PP20[63]);
  UB7_3C63 U98 (W3[65], W8[64], W13[63], PP21[63], PP22[63], PP23[63], PP24[63], PP25[63], PP26[63], PP27[63]);
  UB4_3C63 U99 (W4[65], W9[64], W14[63], PP28[63], PP29[63], PP30[63], PP31[63]);
  UB7_3C64 U100 (W0[66], W5[65], W10[64], PP0[64], PP1[64], PP2[64], PP3[64], PP4[64], PP5[64], PP6[64]);
  UB7_3C64 U101 (W1[66], W6[65], W11[64], PP7[64], PP8[64], PP9[64], PP10[64], PP11[64], PP12[64], PP13[64]);
  UB7_3C64 U102 (W2[66], W7[65], W12[64], PP14[64], PP15[64], PP16[64], PP17[64], PP18[64], PP19[64], PP20[64]);
  UB7_3C64 U103 (W3[66], W8[65], W13[64], PP21[64], PP22[64], PP23[64], PP24[64], PP25[64], PP26[64], PP27[64]);
  UB5_3C64 U104 (W4[66], W9[65], W14[64], PP28[64], PP29[64], PP30[64], PP31[64], PP32[64]);
  UB7_3C65 U105 (W0[67], W5[66], W10[65], PP0[65], PP1[65], PP2[65], PP3[65], PP4[65], PP5[65], PP6[65]);
  UB7_3C65 U106 (W1[67], W6[66], W11[65], PP7[65], PP8[65], PP9[65], PP10[65], PP11[65], PP12[65], PP13[65]);
  UB7_3C65 U107 (W2[67], W7[66], W12[65], PP14[65], PP15[65], PP16[65], PP17[65], PP18[65], PP19[65], PP20[65]);
  UB7_3C65 U108 (W3[67], W8[66], W13[65], PP21[65], PP22[65], PP23[65], PP24[65], PP25[65], PP26[65], PP27[65]);
  UB4_3C65 U109 (W4[67], W9[66], W14[65], PP28[65], PP29[65], PP30[65], PP31[65]);
  UB7_3C66 U110 (W2[68], W5[67], W10[66], PP1[66], PP2[66], PP3[66], PP4[66], PP5[66], PP6[66], PP7[66]);
  UB7_3C66 U111 (W3[68], W6[67], W11[66], PP8[66], PP9[66], PP10[66], PP11[66], PP12[66], PP13[66], PP14[66]);
  UB7_3C66 U112 (W4[68], W7[67], W12[66], PP15[66], PP16[66], PP17[66], PP18[66], PP19[66], PP20[66], PP21[66]);
  UB7_3C66 U113 (W5[68], W8[67], W13[66], PP22[66], PP23[66], PP24[66], PP25[66], PP26[66], PP27[66], PP28[66]);
  UBFA_66 U114 (W9[67], W14[66], PP29[66], PP30[66], PP31[66]);
  UB7_3C67 U115 (W3[69], W6[68], W10[67], PP1[67], PP2[67], PP3[67], PP4[67], PP5[67], PP6[67], PP7[67]);
  UB7_3C67 U116 (W4[69], W7[68], W11[67], PP8[67], PP9[67], PP10[67], PP11[67], PP12[67], PP13[67], PP14[67]);
  UB7_3C67 U117 (W5[69], W8[68], W12[67], PP15[67], PP16[67], PP17[67], PP18[67], PP19[67], PP20[67], PP21[67]);
  UB7_3C67 U118 (W6[69], W9[68], W13[67], PP22[67], PP23[67], PP24[67], PP25[67], PP26[67], PP27[67], PP28[67]);
  UBFA_67 U119 (W10[68], W14[67], PP29[67], PP30[67], PP31[67]);
  UB7_3C68 U120 (W3[70], W7[69], W11[68], PP2[68], PP3[68], PP4[68], PP5[68], PP6[68], PP7[68], PP8[68]);
  UB7_3C68 U121 (W4[70], W8[69], W12[68], PP9[68], PP10[68], PP11[68], PP12[68], PP13[68], PP14[68], PP15[68]);
  UB7_3C68 U122 (W5[70], W9[69], W13[68], PP16[68], PP17[68], PP18[68], PP19[68], PP20[68], PP21[68], PP22[68]);
  UB7_3C68 U123 (W6[70], W10[69], W14[68], PP23[68], PP24[68], PP25[68], PP26[68], PP27[68], PP28[68], PP29[68]);
  UB7_3C69 U124 (W3[71], W7[70], W11[69], PP2[69], PP3[69], PP4[69], PP5[69], PP6[69], PP7[69], PP8[69]);
  UB7_3C69 U125 (W4[71], W8[70], W12[69], PP9[69], PP10[69], PP11[69], PP12[69], PP13[69], PP14[69], PP15[69]);
  UB7_3C69 U126 (W5[71], W9[70], W13[69], PP16[69], PP17[69], PP18[69], PP19[69], PP20[69], PP21[69], PP22[69]);
  UB6_3C69 U127 (W6[71], W10[70], W14[69], PP23[69], PP24[69], PP25[69], PP26[69], PP27[69], PP28[69]);
  UB7_3C70 U128 (W3[72], W7[71], W11[70], PP3[70], PP4[70], PP5[70], PP6[70], PP7[70], PP8[70], PP9[70]);
  UB7_3C70 U129 (W4[72], W8[71], W12[70], PP10[70], PP11[70], PP12[70], PP13[70], PP14[70], PP15[70], PP16[70]);
  UB7_3C70 U130 (W5[72], W9[71], W13[70], PP17[70], PP18[70], PP19[70], PP20[70], PP21[70], PP22[70], PP23[70]);
  UB5_3C70 U131 (W6[72], W10[71], W14[70], PP24[70], PP25[70], PP26[70], PP27[70], PP28[70]);
  UB7_3C71 U132 (W3[73], W7[72], W11[71], PP3[71], PP4[71], PP5[71], PP6[71], PP7[71], PP8[71], PP9[71]);
  UB7_3C71 U133 (W4[73], W8[72], W12[71], PP10[71], PP11[71], PP12[71], PP13[71], PP14[71], PP15[71], PP16[71]);
  UB7_3C71 U134 (W5[73], W9[72], W13[71], PP17[71], PP18[71], PP19[71], PP20[71], PP21[71], PP22[71], PP23[71]);
  UB5_3C71 U135 (W6[73], W10[72], W14[71], PP24[71], PP25[71], PP26[71], PP27[71], PP28[71]);
  UB7_3C72 U136 (W3[74], W7[73], W11[72], PP4[72], PP5[72], PP6[72], PP7[72], PP8[72], PP9[72], PP10[72]);
  UB7_3C72 U137 (W4[74], W8[73], W12[72], PP11[72], PP12[72], PP13[72], PP14[72], PP15[72], PP16[72], PP17[72]);
  UB7_3C72 U138 (W5[74], W9[73], W13[72], PP18[72], PP19[72], PP20[72], PP21[72], PP22[72], PP23[72], PP24[72]);
  UB4_3C72 U139 (W6[74], W10[73], W14[72], PP25[72], PP26[72], PP27[72], PP28[72]);
  UB7_3C73 U140 (W3[75], W7[74], W11[73], PP4[73], PP5[73], PP6[73], PP7[73], PP8[73], PP9[73], PP10[73]);
  UB7_3C73 U141 (W4[75], W8[74], W12[73], PP11[73], PP12[73], PP13[73], PP14[73], PP15[73], PP16[73], PP17[73]);
  UB7_3C73 U142 (W5[75], W9[74], W13[73], PP18[73], PP19[73], PP20[73], PP21[73], PP22[73], PP23[73], PP24[73]);
  UB4_3C73 U143 (W6[75], W10[74], W14[73], PP25[73], PP26[73], PP27[73], PP28[73]);
  UB7_3C74 U144 (W5[76], W7[75], W11[74], PP5[74], PP6[74], PP7[74], PP8[74], PP9[74], PP10[74], PP11[74]);
  UB7_3C74 U145 (W6[76], W8[75], W12[74], PP12[74], PP13[74], PP14[74], PP15[74], PP16[74], PP17[74], PP18[74]);
  UB7_3C74 U146 (W7[76], W9[75], W13[74], PP19[74], PP20[74], PP21[74], PP22[74], PP23[74], PP24[74], PP25[74]);
  UBFA_74 U147 (W10[75], W14[74], PP26[74], PP27[74], PP28[74]);
  UB7_3C75 U148 (W6[77], W8[76], W11[75], PP5[75], PP6[75], PP7[75], PP8[75], PP9[75], PP10[75], PP11[75]);
  UB7_3C75 U149 (W7[77], W9[76], W12[75], PP12[75], PP13[75], PP14[75], PP15[75], PP16[75], PP17[75], PP18[75]);
  UB7_3C75 U150 (W8[77], W10[76], W13[75], PP19[75], PP20[75], PP21[75], PP22[75], PP23[75], PP24[75], PP25[75]);
  UBFA_75 U151 (W11[76], W14[75], PP26[75], PP27[75], PP28[75]);
  UB7_3C76 U152 (W6[78], W9[77], W12[76], PP6[76], PP7[76], PP8[76], PP9[76], PP10[76], PP11[76], PP12[76]);
  UB7_3C76 U153 (W7[78], W10[77], W13[76], PP13[76], PP14[76], PP15[76], PP16[76], PP17[76], PP18[76], PP19[76]);
  UB7_3C76 U154 (W8[78], W11[77], W14[76], PP20[76], PP21[76], PP22[76], PP23[76], PP24[76], PP25[76], PP26[76]);
  UB7_3C77 U155 (W6[79], W9[78], W12[77], PP6[77], PP7[77], PP8[77], PP9[77], PP10[77], PP11[77], PP12[77]);
  UB7_3C77 U156 (W7[79], W10[78], W13[77], PP13[77], PP14[77], PP15[77], PP16[77], PP17[77], PP18[77], PP19[77]);
  UB6_3C77 U157 (W8[79], W11[78], W14[77], PP20[77], PP21[77], PP22[77], PP23[77], PP24[77], PP25[77]);
  UB7_3C78 U158 (W6[80], W9[79], W12[78], PP7[78], PP8[78], PP9[78], PP10[78], PP11[78], PP12[78], PP13[78]);
  UB7_3C78 U159 (W7[80], W10[79], W13[78], PP14[78], PP15[78], PP16[78], PP17[78], PP18[78], PP19[78], PP20[78]);
  UB5_3C78 U160 (W8[80], W11[79], W14[78], PP21[78], PP22[78], PP23[78], PP24[78], PP25[78]);
  UB7_3C79 U161 (W6[81], W9[80], W12[79], PP7[79], PP8[79], PP9[79], PP10[79], PP11[79], PP12[79], PP13[79]);
  UB7_3C79 U162 (W7[81], W10[80], W13[79], PP14[79], PP15[79], PP16[79], PP17[79], PP18[79], PP19[79], PP20[79]);
  UB5_3C79 U163 (W8[81], W11[80], W14[79], PP21[79], PP22[79], PP23[79], PP24[79], PP25[79]);
  UB7_3C80 U164 (W6[82], W9[81], W12[80], PP8[80], PP9[80], PP10[80], PP11[80], PP12[80], PP13[80], PP14[80]);
  UB7_3C80 U165 (W7[82], W10[81], W13[80], PP15[80], PP16[80], PP17[80], PP18[80], PP19[80], PP20[80], PP21[80]);
  UB4_3C80 U166 (W8[82], W11[81], W14[80], PP22[80], PP23[80], PP24[80], PP25[80]);
  UB7_3C81 U167 (W6[83], W9[82], W12[81], PP8[81], PP9[81], PP10[81], PP11[81], PP12[81], PP13[81], PP14[81]);
  UB7_3C81 U168 (W7[83], W10[82], W13[81], PP15[81], PP16[81], PP17[81], PP18[81], PP19[81], PP20[81], PP21[81]);
  UB4_3C81 U169 (W8[83], W11[82], W14[81], PP22[81], PP23[81], PP24[81], PP25[81]);
  UB7_3C82 U170 (W8[84], W9[83], W12[82], PP9[82], PP10[82], PP11[82], PP12[82], PP13[82], PP14[82], PP15[82]);
  UB7_3C82 U171 (W9[84], W10[83], W13[82], PP16[82], PP17[82], PP18[82], PP19[82], PP20[82], PP21[82], PP22[82]);
  UBFA_82 U172 (W11[83], W14[82], PP23[82], PP24[82], PP25[82]);
  UB7_3C83 U173 (W9[85], W10[84], W12[83], PP9[83], PP10[83], PP11[83], PP12[83], PP13[83], PP14[83], PP15[83]);
  UB7_3C83 U174 (W10[85], W11[84], W13[83], PP16[83], PP17[83], PP18[83], PP19[83], PP20[83], PP21[83], PP22[83]);
  UBFA_83 U175 (W12[84], W14[83], PP23[83], PP24[83], PP25[83]);
  UB7_3C84 U176 (W9[86], W11[85], W13[84], PP10[84], PP11[84], PP12[84], PP13[84], PP14[84], PP15[84], PP16[84]);
  UB7_3C84 U177 (W10[86], W12[85], W14[84], PP17[84], PP18[84], PP19[84], PP20[84], PP21[84], PP22[84], PP23[84]);
  UB7_3C85 U178 (W9[87], W11[86], W13[85], PP10[85], PP11[85], PP12[85], PP13[85], PP14[85], PP15[85], PP16[85]);
  UB6_3C85 U179 (W10[87], W12[86], W14[85], PP17[85], PP18[85], PP19[85], PP20[85], PP21[85], PP22[85]);
  UB7_3C86 U180 (W9[88], W11[87], W13[86], PP11[86], PP12[86], PP13[86], PP14[86], PP15[86], PP16[86], PP17[86]);
  UB5_3C86 U181 (W10[88], W12[87], W14[86], PP18[86], PP19[86], PP20[86], PP21[86], PP22[86]);
  UB7_3C87 U182 (W9[89], W11[88], W13[87], PP11[87], PP12[87], PP13[87], PP14[87], PP15[87], PP16[87], PP17[87]);
  UB5_3C87 U183 (W10[89], W12[88], W14[87], PP18[87], PP19[87], PP20[87], PP21[87], PP22[87]);
  UB7_3C88 U184 (W9[90], W11[89], W13[88], PP12[88], PP13[88], PP14[88], PP15[88], PP16[88], PP17[88], PP18[88]);
  UB4_3C88 U185 (W10[90], W12[89], W14[88], PP19[88], PP20[88], PP21[88], PP22[88]);
  UB7_3C89 U186 (W9[91], W11[90], W13[89], PP12[89], PP13[89], PP14[89], PP15[89], PP16[89], PP17[89], PP18[89]);
  UB4_3C89 U187 (W10[91], W12[90], W14[89], PP19[89], PP20[89], PP21[89], PP22[89]);
  UB7_3C90 U188 (W11[92], W11[91], W13[90], PP13[90], PP14[90], PP15[90], PP16[90], PP17[90], PP18[90], PP19[90]);
  UBFA_90 U189 (W12[91], W14[90], PP20[90], PP21[90], PP22[90]);
  UB7_3C91 U190 (W12[93], W12[92], W13[91], PP13[91], PP14[91], PP15[91], PP16[91], PP17[91], PP18[91], PP19[91]);
  UBFA_91 U191 (W13[92], W14[91], PP20[91], PP21[91], PP22[91]);
  UB7_3C92 U192 (W12[94], W13[93], W14[92], PP14[92], PP15[92], PP16[92], PP17[92], PP18[92], PP19[92], PP20[92]);
  UB6_3C93 U193 (W12[95], W13[94], W14[93], PP14[93], PP15[93], PP16[93], PP17[93], PP18[93], PP19[93]);
  UB5_3C94 U194 (W12[96], W13[95], W14[94], PP15[94], PP16[94], PP17[94], PP18[94], PP19[94]);
  UB5_3C95 U195 (W12[97], W13[96], W14[95], PP15[95], PP16[95], PP17[95], PP18[95], PP19[95]);
  UB4_3C96 U196 (W12[98], W13[97], W14[96], PP16[96], PP17[96], PP18[96], PP19[96]);
  UB4_3C97 U197 (W12[99], W13[98], W14[97], PP16[97], PP17[97], PP18[97], PP19[97]);
  UBFA_98 U198 (W13[99], W14[98], PP17[98], PP18[98], PP19[98]);
  UBFA_99 U199 (W14[100], W14[99], PP17[99], PP18[99], PP19[99]);
  UBCON_27_0 U200 (W0[27:0], PP0[27:0]);
  UB1DCON_28 U201 (W0[28], PP2[28]);
  UB1DCON_29 U202 (W0[29], PP3[29]);
  UBCON_31_30 U203 (W0[31:30], PP4[31:30]);
  UBCON_33_32 U204 (W0[33:32], PP6[33:32]);
  UBCON_35_34 U205 (W0[35:34], PP7[35:34]);
  UB1DCON_36 U206 (W0[36], PP9[36]);
  UB1DCON_37 U207 (W0[37], PP10[37]);
  UBCON_39_38 U208 (W0[39:38], PP11[39:38]);
  UBCON_41_40 U209 (W0[41:40], PP13[41:40]);
  UBCON_43_42 U210 (W0[43:42], PP14[43:42]);
  UB1DCON_44 U211 (W0[44], PP16[44]);
  UB1DCON_45 U212 (W0[45], PP17[45]);
  UBCON_47_46 U213 (W0[47:46], PP18[47:46]);
  UBCON_49_48 U214 (W0[49:48], PP20[49:48]);
  UBCON_51_50 U215 (W0[51:50], PP21[51:50]);
  UB1DCON_52 U216 (W0[52], PP23[52]);
  UB1DCON_53 U217 (W0[53], PP24[53]);
  UBCON_55_54 U218 (W0[55:54], PP25[55:54]);
  UBCON_57_56 U219 (W0[57:56], PP27[57:56]);
  UBCON_59_58 U220 (W0[59:58], PP28[59:58]);
  UB1DCON_60 U221 (W0[60], PP30[60]);
  UB1DCON_61 U222 (W0[61], PP31[61]);
  UBCON_63_62 U223 (W0[63:62], PP32[63:62]);
  UB1DCON_68 U224 (W0[68], PP30[68]);
  UBCON_75_69 U225 (W0[75:69], PP29[75:69]);
  UB1DCON_76 U226 (W0[76], PP27[76]);
  UBCON_83_77 U227 (W0[83:77], PP26[83:77]);
  UB1DCON_84 U228 (W0[84], PP24[84]);
  UBCON_91_85 U229 (W0[91:85], PP23[91:85]);
  UB1DCON_92 U230 (W0[92], PP21[92]);
  UBCON_99_93 U231 (W0[99:93], PP20[99:93]);
  UBCON_101_100 U232 (W0[101:100], PP18[101:100]);
  UBCON_103_102 U233 (W0[103:102], PP19[103:102]);
  UBCON_105_104 U234 (W0[105:104], PP20[105:104]);
  UBCON_107_106 U235 (W0[107:106], PP21[107:106]);
  UBCON_109_108 U236 (W0[109:108], PP22[109:108]);
  UBCON_111_110 U237 (W0[111:110], PP23[111:110]);
  UBCON_113_112 U238 (W0[113:112], PP24[113:112]);
  UBCON_115_114 U239 (W0[115:114], PP25[115:114]);
  UBCON_117_116 U240 (W0[117:116], PP26[117:116]);
  UBCON_119_118 U241 (W0[119:118], PP27[119:118]);
  UBCON_121_120 U242 (W0[121:120], PP28[121:120]);
  UBCON_123_122 U243 (W0[123:122], PP29[123:122]);
  UBCON_125_124 U244 (W0[125:124], PP30[125:124]);
  UB1DCON_126 U245 (W0[126], PP31[126]);
  UBCON_27_0 U246 (W1[27:0], PP1[27:0]);
  UB1DCON_28 U247 (W1[28], PP3[28]);
  UB1DCON_29 U248 (W1[29], PP4[29]);
  UBCON_31_30 U249 (W1[31:30], PP5[31:30]);
  UBCON_33_32 U250 (W1[33:32], PP7[33:32]);
  UBCON_35_34 U251 (W1[35:34], PP8[35:34]);
  UB1DCON_36 U252 (W1[36], PP10[36]);
  UB1DCON_37 U253 (W1[37], PP11[37]);
  UBCON_39_38 U254 (W1[39:38], PP12[39:38]);
  UBCON_41_40 U255 (W1[41:40], PP14[41:40]);
  UBCON_43_42 U256 (W1[43:42], PP15[43:42]);
  UB1DCON_44 U257 (W1[44], PP17[44]);
  UB1DCON_45 U258 (W1[45], PP18[45]);
  UBCON_47_46 U259 (W1[47:46], PP19[47:46]);
  UBCON_49_48 U260 (W1[49:48], PP21[49:48]);
  UBCON_51_50 U261 (W1[51:50], PP22[51:50]);
  UB1DCON_52 U262 (W1[52], PP24[52]);
  UB1DCON_53 U263 (W1[53], PP25[53]);
  UBCON_55_54 U264 (W1[55:54], PP26[55:54]);
  UBCON_57_56 U265 (W1[57:56], PP28[57:56]);
  UBCON_59_58 U266 (W1[59:58], PP29[59:58]);
  UB1DCON_60 U267 (W1[60], PP31[60]);
  UB1DCON_68 U268 (W1[68], PP31[68]);
  UBCON_75_69 U269 (W1[75:69], PP30[75:69]);
  UB1DCON_76 U270 (W1[76], PP28[76]);
  UBCON_83_77 U271 (W1[83:77], PP27[83:77]);
  UB1DCON_84 U272 (W1[84], PP25[84]);
  UBCON_91_85 U273 (W1[91:85], PP24[91:85]);
  UB1DCON_92 U274 (W1[92], PP22[92]);
  UBCON_99_93 U275 (W1[99:93], PP21[99:93]);
  UBCON_101_100 U276 (W1[101:100], PP19[101:100]);
  UBCON_103_102 U277 (W1[103:102], PP20[103:102]);
  UBCON_105_104 U278 (W1[105:104], PP21[105:104]);
  UBCON_107_106 U279 (W1[107:106], PP22[107:106]);
  UBCON_109_108 U280 (W1[109:108], PP23[109:108]);
  UBCON_111_110 U281 (W1[111:110], PP24[111:110]);
  UBCON_113_112 U282 (W1[113:112], PP25[113:112]);
  UBCON_115_114 U283 (W1[115:114], PP26[115:114]);
  UBCON_117_116 U284 (W1[117:116], PP27[117:116]);
  UBCON_119_118 U285 (W1[119:118], PP28[119:118]);
  UBCON_121_120 U286 (W1[121:120], PP29[121:120]);
  UBCON_123_122 U287 (W1[123:122], PP30[123:122]);
  UBCON_125_124 U288 (W1[125:124], PP31[125:124]);
  UBCON_27_2 U289 (W2[27:2], PP2[27:2]);
  UB1DCON_28 U290 (W2[28], PP4[28]);
  UB1DCON_29 U291 (W2[29], PP5[29]);
  UBCON_31_30 U292 (W2[31:30], PP6[31:30]);
  UBCON_33_32 U293 (W2[33:32], PP8[33:32]);
  UBCON_35_34 U294 (W2[35:34], PP9[35:34]);
  UB1DCON_36 U295 (W2[36], PP11[36]);
  UB1DCON_37 U296 (W2[37], PP12[37]);
  UBCON_39_38 U297 (W2[39:38], PP13[39:38]);
  UBCON_41_40 U298 (W2[41:40], PP15[41:40]);
  UBCON_43_42 U299 (W2[43:42], PP16[43:42]);
  UB1DCON_44 U300 (W2[44], PP18[44]);
  UB1DCON_45 U301 (W2[45], PP19[45]);
  UBCON_47_46 U302 (W2[47:46], PP20[47:46]);
  UBCON_49_48 U303 (W2[49:48], PP22[49:48]);
  UBCON_51_50 U304 (W2[51:50], PP23[51:50]);
  UB1DCON_52 U305 (W2[52], PP25[52]);
  UB1DCON_53 U306 (W2[53], PP26[53]);
  UBCON_55_54 U307 (W2[55:54], PP27[55:54]);
  UBCON_57_56 U308 (W2[57:56], PP29[57:56]);
  UBCON_59_58 U309 (W2[59:58], PP30[59:58]);
  UBCON_75_69 U310 (W2[75:69], PP31[75:69]);
  UB1DCON_76 U311 (W2[76], PP29[76]);
  UBCON_83_77 U312 (W2[83:77], PP28[83:77]);
  UB1DCON_84 U313 (W2[84], PP26[84]);
  UBCON_91_85 U314 (W2[91:85], PP25[91:85]);
  UB1DCON_92 U315 (W2[92], PP23[92]);
  UBCON_99_93 U316 (W2[99:93], PP22[99:93]);
  UBCON_101_100 U317 (W2[101:100], PP20[101:100]);
  UBCON_103_102 U318 (W2[103:102], PP21[103:102]);
  UBCON_105_104 U319 (W2[105:104], PP22[105:104]);
  UBCON_107_106 U320 (W2[107:106], PP23[107:106]);
  UBCON_109_108 U321 (W2[109:108], PP24[109:108]);
  UBCON_111_110 U322 (W2[111:110], PP25[111:110]);
  UBCON_113_112 U323 (W2[113:112], PP26[113:112]);
  UBCON_115_114 U324 (W2[115:114], PP27[115:114]);
  UBCON_117_116 U325 (W2[117:116], PP28[117:116]);
  UBCON_119_118 U326 (W2[119:118], PP29[119:118]);
  UBCON_121_120 U327 (W2[121:120], PP30[121:120]);
  UBCON_123_122 U328 (W2[123:122], PP31[123:122]);
  UBCON_27_4 U329 (W3[27:4], PP3[27:4]);
  UB1DCON_28 U330 (W3[28], PP5[28]);
  UB1DCON_29 U331 (W3[29], PP6[29]);
  UBCON_31_30 U332 (W3[31:30], PP7[31:30]);
  UBCON_33_32 U333 (W3[33:32], PP9[33:32]);
  UBCON_35_34 U334 (W3[35:34], PP10[35:34]);
  UB1DCON_36 U335 (W3[36], PP12[36]);
  UB1DCON_37 U336 (W3[37], PP13[37]);
  UBCON_39_38 U337 (W3[39:38], PP14[39:38]);
  UBCON_41_40 U338 (W3[41:40], PP16[41:40]);
  UBCON_43_42 U339 (W3[43:42], PP17[43:42]);
  UB1DCON_44 U340 (W3[44], PP19[44]);
  UB1DCON_45 U341 (W3[45], PP20[45]);
  UBCON_47_46 U342 (W3[47:46], PP21[47:46]);
  UBCON_49_48 U343 (W3[49:48], PP23[49:48]);
  UBCON_51_50 U344 (W3[51:50], PP24[51:50]);
  UB1DCON_52 U345 (W3[52], PP26[52]);
  UB1DCON_53 U346 (W3[53], PP27[53]);
  UBCON_55_54 U347 (W3[55:54], PP28[55:54]);
  UB1DCON_76 U348 (W3[76], PP30[76]);
  UBCON_83_77 U349 (W3[83:77], PP29[83:77]);
  UB1DCON_84 U350 (W3[84], PP27[84]);
  UBCON_91_85 U351 (W3[91:85], PP26[91:85]);
  UB1DCON_92 U352 (W3[92], PP24[92]);
  UBCON_99_93 U353 (W3[99:93], PP23[99:93]);
  UBCON_101_100 U354 (W3[101:100], PP21[101:100]);
  UBCON_103_102 U355 (W3[103:102], PP22[103:102]);
  UBCON_105_104 U356 (W3[105:104], PP23[105:104]);
  UBCON_107_106 U357 (W3[107:106], PP24[107:106]);
  UBCON_109_108 U358 (W3[109:108], PP25[109:108]);
  UBCON_111_110 U359 (W3[111:110], PP26[111:110]);
  UBCON_113_112 U360 (W3[113:112], PP27[113:112]);
  UBCON_115_114 U361 (W3[115:114], PP28[115:114]);
  UBCON_117_116 U362 (W3[117:116], PP29[117:116]);
  UBCON_119_118 U363 (W3[119:118], PP30[119:118]);
  UBCON_121_120 U364 (W3[121:120], PP31[121:120]);
  UBCON_27_6 U365 (W4[27:6], PP4[27:6]);
  UB1DCON_28 U366 (W4[28], PP6[28]);
  UB1DCON_29 U367 (W4[29], PP7[29]);
  UBCON_31_30 U368 (W4[31:30], PP8[31:30]);
  UBCON_33_32 U369 (W4[33:32], PP10[33:32]);
  UBCON_35_34 U370 (W4[35:34], PP11[35:34]);
  UB1DCON_36 U371 (W4[36], PP13[36]);
  UB1DCON_37 U372 (W4[37], PP14[37]);
  UBCON_39_38 U373 (W4[39:38], PP15[39:38]);
  UBCON_41_40 U374 (W4[41:40], PP17[41:40]);
  UBCON_43_42 U375 (W4[43:42], PP18[43:42]);
  UB1DCON_44 U376 (W4[44], PP20[44]);
  UB1DCON_45 U377 (W4[45], PP21[45]);
  UBCON_47_46 U378 (W4[47:46], PP22[47:46]);
  UBCON_49_48 U379 (W4[49:48], PP24[49:48]);
  UBCON_51_50 U380 (W4[51:50], PP25[51:50]);
  UB1DCON_52 U381 (W4[52], PP27[52]);
  UB1DCON_76 U382 (W4[76], PP31[76]);
  UBCON_83_77 U383 (W4[83:77], PP30[83:77]);
  UB1DCON_84 U384 (W4[84], PP28[84]);
  UBCON_91_85 U385 (W4[91:85], PP27[91:85]);
  UB1DCON_92 U386 (W4[92], PP25[92]);
  UBCON_99_93 U387 (W4[99:93], PP24[99:93]);
  UBCON_101_100 U388 (W4[101:100], PP22[101:100]);
  UBCON_103_102 U389 (W4[103:102], PP23[103:102]);
  UBCON_105_104 U390 (W4[105:104], PP24[105:104]);
  UBCON_107_106 U391 (W4[107:106], PP25[107:106]);
  UBCON_109_108 U392 (W4[109:108], PP26[109:108]);
  UBCON_111_110 U393 (W4[111:110], PP27[111:110]);
  UBCON_113_112 U394 (W4[113:112], PP28[113:112]);
  UBCON_115_114 U395 (W4[115:114], PP29[115:114]);
  UBCON_117_116 U396 (W4[117:116], PP30[117:116]);
  UBCON_119_118 U397 (W4[119:118], PP31[119:118]);
  UBCON_27_8 U398 (W5[27:8], PP5[27:8]);
  UB1DCON_28 U399 (W5[28], PP7[28]);
  UB1DCON_29 U400 (W5[29], PP8[29]);
  UBCON_31_30 U401 (W5[31:30], PP9[31:30]);
  UBCON_33_32 U402 (W5[33:32], PP11[33:32]);
  UBCON_35_34 U403 (W5[35:34], PP12[35:34]);
  UB1DCON_36 U404 (W5[36], PP14[36]);
  UB1DCON_37 U405 (W5[37], PP15[37]);
  UBCON_39_38 U406 (W5[39:38], PP16[39:38]);
  UBCON_41_40 U407 (W5[41:40], PP18[41:40]);
  UBCON_43_42 U408 (W5[43:42], PP19[43:42]);
  UB1DCON_44 U409 (W5[44], PP21[44]);
  UB1DCON_45 U410 (W5[45], PP22[45]);
  UBCON_47_46 U411 (W5[47:46], PP23[47:46]);
  UBCON_49_48 U412 (W5[49:48], PP25[49:48]);
  UBCON_51_50 U413 (W5[51:50], PP26[51:50]);
  UBCON_83_77 U414 (W5[83:77], PP31[83:77]);
  UB1DCON_84 U415 (W5[84], PP29[84]);
  UBCON_91_85 U416 (W5[91:85], PP28[91:85]);
  UB1DCON_92 U417 (W5[92], PP26[92]);
  UBCON_99_93 U418 (W5[99:93], PP25[99:93]);
  UBCON_101_100 U419 (W5[101:100], PP23[101:100]);
  UBCON_103_102 U420 (W5[103:102], PP24[103:102]);
  UBCON_105_104 U421 (W5[105:104], PP25[105:104]);
  UBCON_107_106 U422 (W5[107:106], PP26[107:106]);
  UBCON_109_108 U423 (W5[109:108], PP27[109:108]);
  UBCON_111_110 U424 (W5[111:110], PP28[111:110]);
  UBCON_113_112 U425 (W5[113:112], PP29[113:112]);
  UBCON_115_114 U426 (W5[115:114], PP30[115:114]);
  UBCON_117_116 U427 (W5[117:116], PP31[117:116]);
  UBCON_27_10 U428 (W6[27:10], PP6[27:10]);
  UB1DCON_28 U429 (W6[28], PP8[28]);
  UB1DCON_29 U430 (W6[29], PP9[29]);
  UBCON_31_30 U431 (W6[31:30], PP10[31:30]);
  UBCON_33_32 U432 (W6[33:32], PP12[33:32]);
  UBCON_35_34 U433 (W6[35:34], PP13[35:34]);
  UB1DCON_36 U434 (W6[36], PP15[36]);
  UB1DCON_37 U435 (W6[37], PP16[37]);
  UBCON_39_38 U436 (W6[39:38], PP17[39:38]);
  UBCON_41_40 U437 (W6[41:40], PP19[41:40]);
  UBCON_43_42 U438 (W6[43:42], PP20[43:42]);
  UB1DCON_44 U439 (W6[44], PP22[44]);
  UB1DCON_45 U440 (W6[45], PP23[45]);
  UBCON_47_46 U441 (W6[47:46], PP24[47:46]);
  UB1DCON_84 U442 (W6[84], PP30[84]);
  UBCON_91_85 U443 (W6[91:85], PP29[91:85]);
  UB1DCON_92 U444 (W6[92], PP27[92]);
  UBCON_99_93 U445 (W6[99:93], PP26[99:93]);
  UBCON_101_100 U446 (W6[101:100], PP24[101:100]);
  UBCON_103_102 U447 (W6[103:102], PP25[103:102]);
  UBCON_105_104 U448 (W6[105:104], PP26[105:104]);
  UBCON_107_106 U449 (W6[107:106], PP27[107:106]);
  UBCON_109_108 U450 (W6[109:108], PP28[109:108]);
  UBCON_111_110 U451 (W6[111:110], PP29[111:110]);
  UBCON_113_112 U452 (W6[113:112], PP30[113:112]);
  UBCON_115_114 U453 (W6[115:114], PP31[115:114]);
  UBCON_27_12 U454 (W7[27:12], PP7[27:12]);
  UB1DCON_28 U455 (W7[28], PP9[28]);
  UB1DCON_29 U456 (W7[29], PP10[29]);
  UBCON_31_30 U457 (W7[31:30], PP11[31:30]);
  UBCON_33_32 U458 (W7[33:32], PP13[33:32]);
  UBCON_35_34 U459 (W7[35:34], PP14[35:34]);
  UB1DCON_36 U460 (W7[36], PP16[36]);
  UB1DCON_37 U461 (W7[37], PP17[37]);
  UBCON_39_38 U462 (W7[39:38], PP18[39:38]);
  UBCON_41_40 U463 (W7[41:40], PP20[41:40]);
  UBCON_43_42 U464 (W7[43:42], PP21[43:42]);
  UB1DCON_44 U465 (W7[44], PP23[44]);
  UB1DCON_84 U466 (W7[84], PP31[84]);
  UBCON_91_85 U467 (W7[91:85], PP30[91:85]);
  UB1DCON_92 U468 (W7[92], PP28[92]);
  UBCON_99_93 U469 (W7[99:93], PP27[99:93]);
  UBCON_101_100 U470 (W7[101:100], PP25[101:100]);
  UBCON_103_102 U471 (W7[103:102], PP26[103:102]);
  UBCON_105_104 U472 (W7[105:104], PP27[105:104]);
  UBCON_107_106 U473 (W7[107:106], PP28[107:106]);
  UBCON_109_108 U474 (W7[109:108], PP29[109:108]);
  UBCON_111_110 U475 (W7[111:110], PP30[111:110]);
  UBCON_113_112 U476 (W7[113:112], PP31[113:112]);
  UBCON_27_14 U477 (W8[27:14], PP8[27:14]);
  UB1DCON_28 U478 (W8[28], PP10[28]);
  UB1DCON_29 U479 (W8[29], PP11[29]);
  UBCON_31_30 U480 (W8[31:30], PP12[31:30]);
  UBCON_33_32 U481 (W8[33:32], PP14[33:32]);
  UBCON_35_34 U482 (W8[35:34], PP15[35:34]);
  UB1DCON_36 U483 (W8[36], PP17[36]);
  UB1DCON_37 U484 (W8[37], PP18[37]);
  UBCON_39_38 U485 (W8[39:38], PP19[39:38]);
  UBCON_41_40 U486 (W8[41:40], PP21[41:40]);
  UBCON_43_42 U487 (W8[43:42], PP22[43:42]);
  UBCON_91_85 U488 (W8[91:85], PP31[91:85]);
  UB1DCON_92 U489 (W8[92], PP29[92]);
  UBCON_99_93 U490 (W8[99:93], PP28[99:93]);
  UBCON_101_100 U491 (W8[101:100], PP26[101:100]);
  UBCON_103_102 U492 (W8[103:102], PP27[103:102]);
  UBCON_105_104 U493 (W8[105:104], PP28[105:104]);
  UBCON_107_106 U494 (W8[107:106], PP29[107:106]);
  UBCON_109_108 U495 (W8[109:108], PP30[109:108]);
  UBCON_111_110 U496 (W8[111:110], PP31[111:110]);
  UBCON_27_16 U497 (W9[27:16], PP9[27:16]);
  UB1DCON_28 U498 (W9[28], PP11[28]);
  UB1DCON_29 U499 (W9[29], PP12[29]);
  UBCON_31_30 U500 (W9[31:30], PP13[31:30]);
  UBCON_33_32 U501 (W9[33:32], PP15[33:32]);
  UBCON_35_34 U502 (W9[35:34], PP16[35:34]);
  UB1DCON_36 U503 (W9[36], PP18[36]);
  UB1DCON_37 U504 (W9[37], PP19[37]);
  UBCON_39_38 U505 (W9[39:38], PP20[39:38]);
  UB1DCON_92 U506 (W9[92], PP30[92]);
  UBCON_99_93 U507 (W9[99:93], PP29[99:93]);
  UBCON_101_100 U508 (W9[101:100], PP27[101:100]);
  UBCON_103_102 U509 (W9[103:102], PP28[103:102]);
  UBCON_105_104 U510 (W9[105:104], PP29[105:104]);
  UBCON_107_106 U511 (W9[107:106], PP30[107:106]);
  UBCON_109_108 U512 (W9[109:108], PP31[109:108]);
  UBCON_27_18 U513 (W10[27:18], PP10[27:18]);
  UB1DCON_28 U514 (W10[28], PP12[28]);
  UB1DCON_29 U515 (W10[29], PP13[29]);
  UBCON_31_30 U516 (W10[31:30], PP14[31:30]);
  UBCON_33_32 U517 (W10[33:32], PP16[33:32]);
  UBCON_35_34 U518 (W10[35:34], PP17[35:34]);
  UB1DCON_36 U519 (W10[36], PP19[36]);
  UB1DCON_92 U520 (W10[92], PP31[92]);
  UBCON_99_93 U521 (W10[99:93], PP30[99:93]);
  UBCON_101_100 U522 (W10[101:100], PP28[101:100]);
  UBCON_103_102 U523 (W10[103:102], PP29[103:102]);
  UBCON_105_104 U524 (W10[105:104], PP30[105:104]);
  UBCON_107_106 U525 (W10[107:106], PP31[107:106]);
  UBCON_27_20 U526 (W11[27:20], PP11[27:20]);
  UB1DCON_28 U527 (W11[28], PP13[28]);
  UB1DCON_29 U528 (W11[29], PP14[29]);
  UBCON_31_30 U529 (W11[31:30], PP15[31:30]);
  UBCON_33_32 U530 (W11[33:32], PP17[33:32]);
  UBCON_35_34 U531 (W11[35:34], PP18[35:34]);
  UBCON_99_93 U532 (W11[99:93], PP31[99:93]);
  UBCON_101_100 U533 (W11[101:100], PP29[101:100]);
  UBCON_103_102 U534 (W11[103:102], PP30[103:102]);
  UBCON_105_104 U535 (W11[105:104], PP31[105:104]);
  UBCON_27_22 U536 (W12[27:22], PP12[27:22]);
  UB1DCON_28 U537 (W12[28], PP14[28]);
  UB1DCON_29 U538 (W12[29], PP15[29]);
  UBCON_31_30 U539 (W12[31:30], PP16[31:30]);
  UBCON_101_100 U540 (W12[101:100], PP30[101:100]);
  UBCON_103_102 U541 (W12[103:102], PP31[103:102]);
  UBCON_27_24 U542 (W13[27:24], PP13[27:24]);
  UB1DCON_28 U543 (W13[28], PP15[28]);
  UBCON_101_100 U544 (W13[101:100], PP31[101:100]);
  UBCON_27_26 U545 (W14[27:26], PP14[27:26]);
  D7_3CTR_126_0_125000 U546 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8, W9, W10, W11, W12, W13, W14);
endmodule

module MultTC_R4B_D73_CS000 (P, IN1, IN2);
  output [127:0] P;
  input [63:0] IN1;
  input [63:0] IN2;
  wire [65:0] PP0;
  wire [67:0] PP1;
  wire [85:18] PP10;
  wire [87:20] PP11;
  wire [89:22] PP12;
  wire [91:24] PP13;
  wire [93:26] PP14;
  wire [95:28] PP15;
  wire [97:30] PP16;
  wire [99:32] PP17;
  wire [101:34] PP18;
  wire [103:36] PP19;
  wire [69:2] PP2;
  wire [105:38] PP20;
  wire [107:40] PP21;
  wire [109:42] PP22;
  wire [111:44] PP23;
  wire [113:46] PP24;
  wire [115:48] PP25;
  wire [117:50] PP26;
  wire [119:52] PP27;
  wire [121:54] PP28;
  wire [123:56] PP29;
  wire [71:4] PP3;
  wire [125:58] PP30;
  wire [126:60] PP31;
  wire [64:62] PP32;
  wire [73:6] PP4;
  wire [75:8] PP5;
  wire [77:10] PP6;
  wire [79:12] PP7;
  wire [81:14] PP8;
  wire [83:16] PP9;
  wire [127:0] P_UB;
  wire [126:0] S1;
  wire [126:0] S2;
  TCR4BPPG_63_0_63_000 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, PP32, IN1, IN2);
  D7_3CTR_65_0_67_0000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, PP32);
  UBCSe_126_0_126_0 U2 (P_UB, S1, S2);
  UBTCCONV127_127_0 U3 (P, P_UB);
endmodule

module TCR4BE_63_0 (O__ds, O__d1, O__d0, I);
  output [31:0] O__ds, O__d1, O__d0;
  input [63:0] I;
  wire [62:0] R;
  wire T;
  TCDECON_63_0 U0 (T, R, I);
  R4BEEL_0_2 U1 (O__ds[0], O__d1[0], O__d0[0], R[1], R[0]);
  R4BEE_1 U2 (O__ds[1], O__d1[1], O__d0[1], R[3], R[2], R[1]);
  R4BEE_2 U3 (O__ds[2], O__d1[2], O__d0[2], R[5], R[4], R[3]);
  R4BEE_3 U4 (O__ds[3], O__d1[3], O__d0[3], R[7], R[6], R[5]);
  R4BEE_4 U5 (O__ds[4], O__d1[4], O__d0[4], R[9], R[8], R[7]);
  R4BEE_5 U6 (O__ds[5], O__d1[5], O__d0[5], R[11], R[10], R[9]);
  R4BEE_6 U7 (O__ds[6], O__d1[6], O__d0[6], R[13], R[12], R[11]);
  R4BEE_7 U8 (O__ds[7], O__d1[7], O__d0[7], R[15], R[14], R[13]);
  R4BEE_8 U9 (O__ds[8], O__d1[8], O__d0[8], R[17], R[16], R[15]);
  R4BEE_9 U10 (O__ds[9], O__d1[9], O__d0[9], R[19], R[18], R[17]);
  R4BEE_10 U11 (O__ds[10], O__d1[10], O__d0[10], R[21], R[20], R[19]);
  R4BEE_11 U12 (O__ds[11], O__d1[11], O__d0[11], R[23], R[22], R[21]);
  R4BEE_12 U13 (O__ds[12], O__d1[12], O__d0[12], R[25], R[24], R[23]);
  R4BEE_13 U14 (O__ds[13], O__d1[13], O__d0[13], R[27], R[26], R[25]);
  R4BEE_14 U15 (O__ds[14], O__d1[14], O__d0[14], R[29], R[28], R[27]);
  R4BEE_15 U16 (O__ds[15], O__d1[15], O__d0[15], R[31], R[30], R[29]);
  R4BEE_16 U17 (O__ds[16], O__d1[16], O__d0[16], R[33], R[32], R[31]);
  R4BEE_17 U18 (O__ds[17], O__d1[17], O__d0[17], R[35], R[34], R[33]);
  R4BEE_18 U19 (O__ds[18], O__d1[18], O__d0[18], R[37], R[36], R[35]);
  R4BEE_19 U20 (O__ds[19], O__d1[19], O__d0[19], R[39], R[38], R[37]);
  R4BEE_20 U21 (O__ds[20], O__d1[20], O__d0[20], R[41], R[40], R[39]);
  R4BEE_21 U22 (O__ds[21], O__d1[21], O__d0[21], R[43], R[42], R[41]);
  R4BEE_22 U23 (O__ds[22], O__d1[22], O__d0[22], R[45], R[44], R[43]);
  R4BEE_23 U24 (O__ds[23], O__d1[23], O__d0[23], R[47], R[46], R[45]);
  R4BEE_24 U25 (O__ds[24], O__d1[24], O__d0[24], R[49], R[48], R[47]);
  R4BEE_25 U26 (O__ds[25], O__d1[25], O__d0[25], R[51], R[50], R[49]);
  R4BEE_26 U27 (O__ds[26], O__d1[26], O__d0[26], R[53], R[52], R[51]);
  R4BEE_27 U28 (O__ds[27], O__d1[27], O__d0[27], R[55], R[54], R[53]);
  R4BEE_28 U29 (O__ds[28], O__d1[28], O__d0[28], R[57], R[56], R[55]);
  R4BEE_29 U30 (O__ds[29], O__d1[29], O__d0[29], R[59], R[58], R[57]);
  R4BEE_30 U31 (O__ds[30], O__d1[30], O__d0[30], R[61], R[60], R[59]);
  R4BEEH_31_3 U32 (O__ds[31], O__d1[31], O__d0[31], T, R[62], R[61]);
endmodule

module TCR4BPPG_63_0_63_000 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, PP32, IN1, IN2);
  output [65:0] PP0;
  output [67:0] PP1;
  output [85:18] PP10;
  output [87:20] PP11;
  output [89:22] PP12;
  output [91:24] PP13;
  output [93:26] PP14;
  output [95:28] PP15;
  output [97:30] PP16;
  output [99:32] PP17;
  output [101:34] PP18;
  output [103:36] PP19;
  output [69:2] PP2;
  output [105:38] PP20;
  output [107:40] PP21;
  output [109:42] PP22;
  output [111:44] PP23;
  output [113:46] PP24;
  output [115:48] PP25;
  output [117:50] PP26;
  output [119:52] PP27;
  output [121:54] PP28;
  output [123:56] PP29;
  output [71:4] PP3;
  output [125:58] PP30;
  output [126:60] PP31;
  output [64:62] PP32;
  output [73:6] PP4;
  output [75:8] PP5;
  output [77:10] PP6;
  output [79:12] PP7;
  output [81:14] PP8;
  output [83:16] PP9;
  input [63:0] IN1;
  input [63:0] IN2;
  wire B0;
  wire B1;
  wire B10;
  wire B11;
  wire B12;
  wire B13;
  wire B14;
  wire B15;
  wire B16;
  wire B17;
  wire B18;
  wire B19;
  wire B2;
  wire B20;
  wire B21;
  wire B22;
  wire B23;
  wire B24;
  wire B25;
  wire B26;
  wire B27;
  wire B28;
  wire B29;
  wire B3;
  wire B30;
  wire B31;
  wire B4;
  wire B5;
  wire B6;
  wire B7;
  wire B8;
  wire B9;
  wire [31:0] IN2SD__ds, IN2SD__d1, IN2SD__d0;
  wire [64:0] PPT0;
  wire [66:2] PPT1;
  wire [84:20] PPT10;
  wire [86:22] PPT11;
  wire [88:24] PPT12;
  wire [90:26] PPT13;
  wire [92:28] PPT14;
  wire [94:30] PPT15;
  wire [96:32] PPT16;
  wire [98:34] PPT17;
  wire [100:36] PPT18;
  wire [102:38] PPT19;
  wire [68:4] PPT2;
  wire [104:40] PPT20;
  wire [106:42] PPT21;
  wire [108:44] PPT22;
  wire [110:46] PPT23;
  wire [112:48] PPT24;
  wire [114:50] PPT25;
  wire [116:52] PPT26;
  wire [118:54] PPT27;
  wire [120:56] PPT28;
  wire [122:58] PPT29;
  wire [70:6] PPT3;
  wire [124:60] PPT30;
  wire [126:62] PPT31;
  wire [72:8] PPT4;
  wire [74:10] PPT5;
  wire [76:12] PPT6;
  wire [78:14] PPT7;
  wire [80:16] PPT8;
  wire [82:18] PPT9;
  wire S0;
  wire S1;
  wire S10;
  wire S11;
  wire S12;
  wire S13;
  wire S14;
  wire S15;
  wire S16;
  wire S17;
  wire S18;
  wire S19;
  wire S2;
  wire S20;
  wire S21;
  wire S22;
  wire S23;
  wire S24;
  wire S25;
  wire S26;
  wire S27;
  wire S28;
  wire S29;
  wire S3;
  wire S30;
  wire S31;
  wire S4;
  wire S5;
  wire S6;
  wire S7;
  wire S8;
  wire S9;
  TCR4BE_63_0 U0 (IN2SD__ds, IN2SD__d1, IN2SD__d0, IN2);
  TCSD4VPPG_63_0_0 U1 (PPT0, S0, IN1, IN2SD__ds[0], IN2SD__d1[0], IN2SD__d0[0]);
  TCSD4VPPG_63_0_1 U2 (PPT1, S1, IN1, IN2SD__ds[1], IN2SD__d1[1], IN2SD__d0[1]);
  TCSD4VPPG_63_0_2 U3 (PPT2, S2, IN1, IN2SD__ds[2], IN2SD__d1[2], IN2SD__d0[2]);
  TCSD4VPPG_63_0_3 U4 (PPT3, S3, IN1, IN2SD__ds[3], IN2SD__d1[3], IN2SD__d0[3]);
  TCSD4VPPG_63_0_4 U5 (PPT4, S4, IN1, IN2SD__ds[4], IN2SD__d1[4], IN2SD__d0[4]);
  TCSD4VPPG_63_0_5 U6 (PPT5, S5, IN1, IN2SD__ds[5], IN2SD__d1[5], IN2SD__d0[5]);
  TCSD4VPPG_63_0_6 U7 (PPT6, S6, IN1, IN2SD__ds[6], IN2SD__d1[6], IN2SD__d0[6]);
  TCSD4VPPG_63_0_7 U8 (PPT7, S7, IN1, IN2SD__ds[7], IN2SD__d1[7], IN2SD__d0[7]);
  TCSD4VPPG_63_0_8 U9 (PPT8, S8, IN1, IN2SD__ds[8], IN2SD__d1[8], IN2SD__d0[8]);
  TCSD4VPPG_63_0_9 U10 (PPT9, S9, IN1, IN2SD__ds[9], IN2SD__d1[9], IN2SD__d0[9]);
  TCSD4VPPG_63_0_10 U11 (PPT10, S10, IN1, IN2SD__ds[10], IN2SD__d1[10], IN2SD__d0[10]);
  TCSD4VPPG_63_0_11 U12 (PPT11, S11, IN1, IN2SD__ds[11], IN2SD__d1[11], IN2SD__d0[11]);
  TCSD4VPPG_63_0_12 U13 (PPT12, S12, IN1, IN2SD__ds[12], IN2SD__d1[12], IN2SD__d0[12]);
  TCSD4VPPG_63_0_13 U14 (PPT13, S13, IN1, IN2SD__ds[13], IN2SD__d1[13], IN2SD__d0[13]);
  TCSD4VPPG_63_0_14 U15 (PPT14, S14, IN1, IN2SD__ds[14], IN2SD__d1[14], IN2SD__d0[14]);
  TCSD4VPPG_63_0_15 U16 (PPT15, S15, IN1, IN2SD__ds[15], IN2SD__d1[15], IN2SD__d0[15]);
  TCSD4VPPG_63_0_16 U17 (PPT16, S16, IN1, IN2SD__ds[16], IN2SD__d1[16], IN2SD__d0[16]);
  TCSD4VPPG_63_0_17 U18 (PPT17, S17, IN1, IN2SD__ds[17], IN2SD__d1[17], IN2SD__d0[17]);
  TCSD4VPPG_63_0_18 U19 (PPT18, S18, IN1, IN2SD__ds[18], IN2SD__d1[18], IN2SD__d0[18]);
  TCSD4VPPG_63_0_19 U20 (PPT19, S19, IN1, IN2SD__ds[19], IN2SD__d1[19], IN2SD__d0[19]);
  TCSD4VPPG_63_0_20 U21 (PPT20, S20, IN1, IN2SD__ds[20], IN2SD__d1[20], IN2SD__d0[20]);
  TCSD4VPPG_63_0_21 U22 (PPT21, S21, IN1, IN2SD__ds[21], IN2SD__d1[21], IN2SD__d0[21]);
  TCSD4VPPG_63_0_22 U23 (PPT22, S22, IN1, IN2SD__ds[22], IN2SD__d1[22], IN2SD__d0[22]);
  TCSD4VPPG_63_0_23 U24 (PPT23, S23, IN1, IN2SD__ds[23], IN2SD__d1[23], IN2SD__d0[23]);
  TCSD4VPPG_63_0_24 U25 (PPT24, S24, IN1, IN2SD__ds[24], IN2SD__d1[24], IN2SD__d0[24]);
  TCSD4VPPG_63_0_25 U26 (PPT25, S25, IN1, IN2SD__ds[25], IN2SD__d1[25], IN2SD__d0[25]);
  TCSD4VPPG_63_0_26 U27 (PPT26, S26, IN1, IN2SD__ds[26], IN2SD__d1[26], IN2SD__d0[26]);
  TCSD4VPPG_63_0_27 U28 (PPT27, S27, IN1, IN2SD__ds[27], IN2SD__d1[27], IN2SD__d0[27]);
  TCSD4VPPG_63_0_28 U29 (PPT28, S28, IN1, IN2SD__ds[28], IN2SD__d1[28], IN2SD__d0[28]);
  TCSD4VPPG_63_0_29 U30 (PPT29, S29, IN1, IN2SD__ds[29], IN2SD__d1[29], IN2SD__d0[29]);
  TCSD4VPPG_63_0_30 U31 (PPT30, S30, IN1, IN2SD__ds[30], IN2SD__d1[30], IN2SD__d0[30]);
  TCSD4VPPG_63_0_31 U32 (PPT31, S31, IN1, IN2SD__ds[31], IN2SD__d1[31], IN2SD__d0[31]);
  UBOne_65 U33 (B0);
  UBCMBIN_65_65_64_000 U34 (PP0, B0, PPT0);
  UBOne_67 U35 (B1);
  UBCMBIN_67_67_66_000 U36 (PP1, B1, PPT1, S0);
  UBOne_69 U37 (B2);
  UBCMBIN_69_69_68_000 U38 (PP2, B2, PPT2, S1);
  UBOne_71 U39 (B3);
  UBCMBIN_71_71_70_000 U40 (PP3, B3, PPT3, S2);
  UBOne_73 U41 (B4);
  UBCMBIN_73_73_72_000 U42 (PP4, B4, PPT4, S3);
  UBOne_75 U43 (B5);
  UBCMBIN_75_75_74_000 U44 (PP5, B5, PPT5, S4);
  UBOne_77 U45 (B6);
  UBCMBIN_77_77_76_000 U46 (PP6, B6, PPT6, S5);
  UBOne_79 U47 (B7);
  UBCMBIN_79_79_78_000 U48 (PP7, B7, PPT7, S6);
  UBOne_81 U49 (B8);
  UBCMBIN_81_81_80_000 U50 (PP8, B8, PPT8, S7);
  UBOne_83 U51 (B9);
  UBCMBIN_83_83_82_000 U52 (PP9, B9, PPT9, S8);
  UBOne_85 U53 (B10);
  UBCMBIN_85_85_84_000 U54 (PP10, B10, PPT10, S9);
  UBOne_87 U55 (B11);
  UBCMBIN_87_87_86_000 U56 (PP11, B11, PPT11, S10);
  UBOne_89 U57 (B12);
  UBCMBIN_89_89_88_000 U58 (PP12, B12, PPT12, S11);
  UBOne_91 U59 (B13);
  UBCMBIN_91_91_90_000 U60 (PP13, B13, PPT13, S12);
  UBOne_93 U61 (B14);
  UBCMBIN_93_93_92_000 U62 (PP14, B14, PPT14, S13);
  UBOne_95 U63 (B15);
  UBCMBIN_95_95_94_000 U64 (PP15, B15, PPT15, S14);
  UBOne_97 U65 (B16);
  UBCMBIN_97_97_96_000 U66 (PP16, B16, PPT16, S15);
  UBOne_99 U67 (B17);
  UBCMBIN_99_99_98_000 U68 (PP17, B17, PPT17, S16);
  UBOne_101 U69 (B18);
  UBCMBIN_101_101_1000 U70 (PP18, B18, PPT18, S17);
  UBOne_103 U71 (B19);
  UBCMBIN_103_103_1000 U72 (PP19, B19, PPT19, S18);
  UBOne_105 U73 (B20);
  UBCMBIN_105_105_1000 U74 (PP20, B20, PPT20, S19);
  UBOne_107 U75 (B21);
  UBCMBIN_107_107_1000 U76 (PP21, B21, PPT21, S20);
  UBOne_109 U77 (B22);
  UBCMBIN_109_109_1000 U78 (PP22, B22, PPT22, S21);
  UBOne_111 U79 (B23);
  UBCMBIN_111_111_1000 U80 (PP23, B23, PPT23, S22);
  UBOne_113 U81 (B24);
  UBCMBIN_113_113_1000 U82 (PP24, B24, PPT24, S23);
  UBOne_115 U83 (B25);
  UBCMBIN_115_115_1000 U84 (PP25, B25, PPT25, S24);
  UBOne_117 U85 (B26);
  UBCMBIN_117_117_1000 U86 (PP26, B26, PPT26, S25);
  UBOne_119 U87 (B27);
  UBCMBIN_119_119_1000 U88 (PP27, B27, PPT27, S26);
  UBOne_121 U89 (B28);
  UBCMBIN_121_121_1000 U90 (PP28, B28, PPT28, S27);
  UBOne_123 U91 (B29);
  UBCMBIN_123_123_1000 U92 (PP29, B29, PPT29, S28);
  UBOne_125 U93 (B30);
  UBCMBIN_125_125_1000 U94 (PP30, B30, PPT30, S29);
  UBCMBIN_126_62_60000 U95 (PP31, PPT31, S30);
  UBOne_64 U96 (B31);
  UBCMBIN_64_64_62_000 U97 (PP32, B31, S31);
endmodule

module TCSD4VPPG_63_0_0 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [64:0] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [63:0] W_R;
  wire W_T;
  SD41DDECON_0 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_0 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_64_0 U3 (PP, W_T, W_R, S);
  UBBBG_0 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_1 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [66:2] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [65:2] W_R;
  wire W_T;
  SD41DDECON_1 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_1 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_66_2 U3 (PP, W_T, W_R, S);
  UBBBG_2 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_10 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [84:20] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [83:20] W_R;
  wire W_T;
  SD41DDECON_10 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_10 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_84_20 U3 (PP, W_T, W_R, S);
  UBBBG_20 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_11 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [86:22] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [85:22] W_R;
  wire W_T;
  SD41DDECON_11 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_11 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_86_22 U3 (PP, W_T, W_R, S);
  UBBBG_22 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_12 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [88:24] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [87:24] W_R;
  wire W_T;
  SD41DDECON_12 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_12 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_88_24 U3 (PP, W_T, W_R, S);
  UBBBG_24 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_13 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [90:26] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [89:26] W_R;
  wire W_T;
  SD41DDECON_13 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_13 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_90_26 U3 (PP, W_T, W_R, S);
  UBBBG_26 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_14 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [92:28] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [91:28] W_R;
  wire W_T;
  SD41DDECON_14 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_14 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_92_28 U3 (PP, W_T, W_R, S);
  UBBBG_28 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_15 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [94:30] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [93:30] W_R;
  wire W_T;
  SD41DDECON_15 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_15 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_94_30 U3 (PP, W_T, W_R, S);
  UBBBG_30 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_16 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [96:32] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [95:32] W_R;
  wire W_T;
  SD41DDECON_16 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_16 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_96_32 U3 (PP, W_T, W_R, S);
  UBBBG_32 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_17 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [98:34] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [97:34] W_R;
  wire W_T;
  SD41DDECON_17 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_17 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_98_34 U3 (PP, W_T, W_R, S);
  UBBBG_34 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_18 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [100:36] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [99:36] W_R;
  wire W_T;
  SD41DDECON_18 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_18 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_100_36 U3 (PP, W_T, W_R, S);
  UBBBG_36 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_19 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [102:38] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [101:38] W_R;
  wire W_T;
  SD41DDECON_19 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_19 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_102_38 U3 (PP, W_T, W_R, S);
  UBBBG_38 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_2 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [68:4] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [67:4] W_R;
  wire W_T;
  SD41DDECON_2 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_2 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_68_4 U3 (PP, W_T, W_R, S);
  UBBBG_4 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_20 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [104:40] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [103:40] W_R;
  wire W_T;
  SD41DDECON_20 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_20 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_104_40 U3 (PP, W_T, W_R, S);
  UBBBG_40 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_21 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [106:42] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [105:42] W_R;
  wire W_T;
  SD41DDECON_21 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_21 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_106_42 U3 (PP, W_T, W_R, S);
  UBBBG_42 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_22 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [108:44] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [107:44] W_R;
  wire W_T;
  SD41DDECON_22 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_22 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_108_44 U3 (PP, W_T, W_R, S);
  UBBBG_44 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_23 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [110:46] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [109:46] W_R;
  wire W_T;
  SD41DDECON_23 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_23 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_110_46 U3 (PP, W_T, W_R, S);
  UBBBG_46 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_24 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [112:48] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [111:48] W_R;
  wire W_T;
  SD41DDECON_24 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_24 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_112_48 U3 (PP, W_T, W_R, S);
  UBBBG_48 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_25 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [114:50] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [113:50] W_R;
  wire W_T;
  SD41DDECON_25 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_25 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_114_50 U3 (PP, W_T, W_R, S);
  UBBBG_50 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_26 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [116:52] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [115:52] W_R;
  wire W_T;
  SD41DDECON_26 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_26 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_116_52 U3 (PP, W_T, W_R, S);
  UBBBG_52 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_27 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [118:54] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [117:54] W_R;
  wire W_T;
  SD41DDECON_27 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_27 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_118_54 U3 (PP, W_T, W_R, S);
  UBBBG_54 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_28 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [120:56] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [119:56] W_R;
  wire W_T;
  SD41DDECON_28 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_28 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_120_56 U3 (PP, W_T, W_R, S);
  UBBBG_56 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_29 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [122:58] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [121:58] W_R;
  wire W_T;
  SD41DDECON_29 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_29 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_122_58 U3 (PP, W_T, W_R, S);
  UBBBG_58 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_3 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [70:6] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [69:6] W_R;
  wire W_T;
  SD41DDECON_3 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_3 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_70_6 U3 (PP, W_T, W_R, S);
  UBBBG_6 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_30 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [124:60] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [123:60] W_R;
  wire W_T;
  SD41DDECON_30 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_30 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_124_60 U3 (PP, W_T, W_R, S);
  UBBBG_60 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_31 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [126:62] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [125:62] W_R;
  wire W_T;
  SD41DDECON_31 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_31 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_126_62 U3 (PP, W_T, W_R, S);
  UBBBG_62 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_4 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [72:8] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [71:8] W_R;
  wire W_T;
  SD41DDECON_4 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_4 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_72_8 U3 (PP, W_T, W_R, S);
  UBBBG_8 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_5 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [74:10] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [73:10] W_R;
  wire W_T;
  SD41DDECON_5 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_5 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_74_10 U3 (PP, W_T, W_R, S);
  UBBBG_10 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_6 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [76:12] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [75:12] W_R;
  wire W_T;
  SD41DDECON_6 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_6 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_76_12 U3 (PP, W_T, W_R, S);
  UBBBG_12 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_7 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [78:14] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [77:14] W_R;
  wire W_T;
  SD41DDECON_7 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_7 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_78_14 U3 (PP, W_T, W_R, S);
  UBBBG_14 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_8 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [80:16] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [79:16] W_R;
  wire W_T;
  SD41DDECON_8 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_8 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_80_16 U3 (PP, W_T, W_R, S);
  UBBBG_16 U4 (C, S);
endmodule

module TCSD4VPPG_63_0_9 (PP, C, IN1, IN2__ds, IN2__d1, IN2__d0);
  output C;
  output [82:18] PP;
  input [63:0] IN1;
  input IN2__ds, IN2__d1, IN2__d0;
  wire [62:0] IN1_R;
  wire IN1_T;
  wire S;
  wire U__d1, U__d0;
  wire [81:18] W_R;
  wire W_T;
  SD41DDECON_9 U0 (S, U__d1, U__d0, IN2__ds, IN2__d1, IN2__d0);
  TCDECON_63_0 U1 (IN1_T, IN1_R, IN1);
  TCU4VPPG_63_0_9 U2 (W_T, W_R, IN1_T, IN1_R, U__d1, U__d0);
  TUBWCON_82_18 U3 (PP, W_T, W_R, S);
  UBBBG_18 U4 (C, S);
endmodule

module TCU4VPPG_63_0_0 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [63:0] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [63:1] P;
  U4DPPGL_0_0 U0 (P[1], O_R[0], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_0 U1 (P[2], O_R[1], IN1_R[1], U__d1, U__d0, P[1]);
  U4DPPG_2_0 U2 (P[3], O_R[2], IN1_R[2], U__d1, U__d0, P[2]);
  U4DPPG_3_0 U3 (P[4], O_R[3], IN1_R[3], U__d1, U__d0, P[3]);
  U4DPPG_4_0 U4 (P[5], O_R[4], IN1_R[4], U__d1, U__d0, P[4]);
  U4DPPG_5_0 U5 (P[6], O_R[5], IN1_R[5], U__d1, U__d0, P[5]);
  U4DPPG_6_0 U6 (P[7], O_R[6], IN1_R[6], U__d1, U__d0, P[6]);
  U4DPPG_7_0 U7 (P[8], O_R[7], IN1_R[7], U__d1, U__d0, P[7]);
  U4DPPG_8_0 U8 (P[9], O_R[8], IN1_R[8], U__d1, U__d0, P[8]);
  U4DPPG_9_0 U9 (P[10], O_R[9], IN1_R[9], U__d1, U__d0, P[9]);
  U4DPPG_10_0 U10 (P[11], O_R[10], IN1_R[10], U__d1, U__d0, P[10]);
  U4DPPG_11_0 U11 (P[12], O_R[11], IN1_R[11], U__d1, U__d0, P[11]);
  U4DPPG_12_0 U12 (P[13], O_R[12], IN1_R[12], U__d1, U__d0, P[12]);
  U4DPPG_13_0 U13 (P[14], O_R[13], IN1_R[13], U__d1, U__d0, P[13]);
  U4DPPG_14_0 U14 (P[15], O_R[14], IN1_R[14], U__d1, U__d0, P[14]);
  U4DPPG_15_0 U15 (P[16], O_R[15], IN1_R[15], U__d1, U__d0, P[15]);
  U4DPPG_16_0 U16 (P[17], O_R[16], IN1_R[16], U__d1, U__d0, P[16]);
  U4DPPG_17_0 U17 (P[18], O_R[17], IN1_R[17], U__d1, U__d0, P[17]);
  U4DPPG_18_0 U18 (P[19], O_R[18], IN1_R[18], U__d1, U__d0, P[18]);
  U4DPPG_19_0 U19 (P[20], O_R[19], IN1_R[19], U__d1, U__d0, P[19]);
  U4DPPG_20_0 U20 (P[21], O_R[20], IN1_R[20], U__d1, U__d0, P[20]);
  U4DPPG_21_0 U21 (P[22], O_R[21], IN1_R[21], U__d1, U__d0, P[21]);
  U4DPPG_22_0 U22 (P[23], O_R[22], IN1_R[22], U__d1, U__d0, P[22]);
  U4DPPG_23_0 U23 (P[24], O_R[23], IN1_R[23], U__d1, U__d0, P[23]);
  U4DPPG_24_0 U24 (P[25], O_R[24], IN1_R[24], U__d1, U__d0, P[24]);
  U4DPPG_25_0 U25 (P[26], O_R[25], IN1_R[25], U__d1, U__d0, P[25]);
  U4DPPG_26_0 U26 (P[27], O_R[26], IN1_R[26], U__d1, U__d0, P[26]);
  U4DPPG_27_0 U27 (P[28], O_R[27], IN1_R[27], U__d1, U__d0, P[27]);
  U4DPPG_28_0 U28 (P[29], O_R[28], IN1_R[28], U__d1, U__d0, P[28]);
  U4DPPG_29_0 U29 (P[30], O_R[29], IN1_R[29], U__d1, U__d0, P[29]);
  U4DPPG_30_0 U30 (P[31], O_R[30], IN1_R[30], U__d1, U__d0, P[30]);
  U4DPPG_31_0 U31 (P[32], O_R[31], IN1_R[31], U__d1, U__d0, P[31]);
  U4DPPG_32_0 U32 (P[33], O_R[32], IN1_R[32], U__d1, U__d0, P[32]);
  U4DPPG_33_0 U33 (P[34], O_R[33], IN1_R[33], U__d1, U__d0, P[33]);
  U4DPPG_34_0 U34 (P[35], O_R[34], IN1_R[34], U__d1, U__d0, P[34]);
  U4DPPG_35_0 U35 (P[36], O_R[35], IN1_R[35], U__d1, U__d0, P[35]);
  U4DPPG_36_0 U36 (P[37], O_R[36], IN1_R[36], U__d1, U__d0, P[36]);
  U4DPPG_37_0 U37 (P[38], O_R[37], IN1_R[37], U__d1, U__d0, P[37]);
  U4DPPG_38_0 U38 (P[39], O_R[38], IN1_R[38], U__d1, U__d0, P[38]);
  U4DPPG_39_0 U39 (P[40], O_R[39], IN1_R[39], U__d1, U__d0, P[39]);
  U4DPPG_40_0 U40 (P[41], O_R[40], IN1_R[40], U__d1, U__d0, P[40]);
  U4DPPG_41_0 U41 (P[42], O_R[41], IN1_R[41], U__d1, U__d0, P[41]);
  U4DPPG_42_0 U42 (P[43], O_R[42], IN1_R[42], U__d1, U__d0, P[42]);
  U4DPPG_43_0 U43 (P[44], O_R[43], IN1_R[43], U__d1, U__d0, P[43]);
  U4DPPG_44_0 U44 (P[45], O_R[44], IN1_R[44], U__d1, U__d0, P[44]);
  U4DPPG_45_0 U45 (P[46], O_R[45], IN1_R[45], U__d1, U__d0, P[45]);
  U4DPPG_46_0 U46 (P[47], O_R[46], IN1_R[46], U__d1, U__d0, P[46]);
  U4DPPG_47_0 U47 (P[48], O_R[47], IN1_R[47], U__d1, U__d0, P[47]);
  U4DPPG_48_0 U48 (P[49], O_R[48], IN1_R[48], U__d1, U__d0, P[48]);
  U4DPPG_49_0 U49 (P[50], O_R[49], IN1_R[49], U__d1, U__d0, P[49]);
  U4DPPG_50_0 U50 (P[51], O_R[50], IN1_R[50], U__d1, U__d0, P[50]);
  U4DPPG_51_0 U51 (P[52], O_R[51], IN1_R[51], U__d1, U__d0, P[51]);
  U4DPPG_52_0 U52 (P[53], O_R[52], IN1_R[52], U__d1, U__d0, P[52]);
  U4DPPG_53_0 U53 (P[54], O_R[53], IN1_R[53], U__d1, U__d0, P[53]);
  U4DPPG_54_0 U54 (P[55], O_R[54], IN1_R[54], U__d1, U__d0, P[54]);
  U4DPPG_55_0 U55 (P[56], O_R[55], IN1_R[55], U__d1, U__d0, P[55]);
  U4DPPG_56_0 U56 (P[57], O_R[56], IN1_R[56], U__d1, U__d0, P[56]);
  U4DPPG_57_0 U57 (P[58], O_R[57], IN1_R[57], U__d1, U__d0, P[57]);
  U4DPPG_58_0 U58 (P[59], O_R[58], IN1_R[58], U__d1, U__d0, P[58]);
  U4DPPG_59_0 U59 (P[60], O_R[59], IN1_R[59], U__d1, U__d0, P[59]);
  U4DPPG_60_0 U60 (P[61], O_R[60], IN1_R[60], U__d1, U__d0, P[60]);
  U4DPPG_61_0 U61 (P[62], O_R[61], IN1_R[61], U__d1, U__d0, P[61]);
  U4DPPG_62_0 U62 (P[63], O_R[62], IN1_R[62], U__d1, U__d0, P[62]);
  U4DPPGH_63_0 U63 (O_T, O_R[63], IN1_T, U__d1, U__d0, P[63]);
endmodule

module TCU4VPPG_63_0_1 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [65:2] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [65:3] P;
  U4DPPGL_0_1 U0 (P[3], O_R[2], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_1 U1 (P[4], O_R[3], IN1_R[1], U__d1, U__d0, P[3]);
  U4DPPG_2_1 U2 (P[5], O_R[4], IN1_R[2], U__d1, U__d0, P[4]);
  U4DPPG_3_1 U3 (P[6], O_R[5], IN1_R[3], U__d1, U__d0, P[5]);
  U4DPPG_4_1 U4 (P[7], O_R[6], IN1_R[4], U__d1, U__d0, P[6]);
  U4DPPG_5_1 U5 (P[8], O_R[7], IN1_R[5], U__d1, U__d0, P[7]);
  U4DPPG_6_1 U6 (P[9], O_R[8], IN1_R[6], U__d1, U__d0, P[8]);
  U4DPPG_7_1 U7 (P[10], O_R[9], IN1_R[7], U__d1, U__d0, P[9]);
  U4DPPG_8_1 U8 (P[11], O_R[10], IN1_R[8], U__d1, U__d0, P[10]);
  U4DPPG_9_1 U9 (P[12], O_R[11], IN1_R[9], U__d1, U__d0, P[11]);
  U4DPPG_10_1 U10 (P[13], O_R[12], IN1_R[10], U__d1, U__d0, P[12]);
  U4DPPG_11_1 U11 (P[14], O_R[13], IN1_R[11], U__d1, U__d0, P[13]);
  U4DPPG_12_1 U12 (P[15], O_R[14], IN1_R[12], U__d1, U__d0, P[14]);
  U4DPPG_13_1 U13 (P[16], O_R[15], IN1_R[13], U__d1, U__d0, P[15]);
  U4DPPG_14_1 U14 (P[17], O_R[16], IN1_R[14], U__d1, U__d0, P[16]);
  U4DPPG_15_1 U15 (P[18], O_R[17], IN1_R[15], U__d1, U__d0, P[17]);
  U4DPPG_16_1 U16 (P[19], O_R[18], IN1_R[16], U__d1, U__d0, P[18]);
  U4DPPG_17_1 U17 (P[20], O_R[19], IN1_R[17], U__d1, U__d0, P[19]);
  U4DPPG_18_1 U18 (P[21], O_R[20], IN1_R[18], U__d1, U__d0, P[20]);
  U4DPPG_19_1 U19 (P[22], O_R[21], IN1_R[19], U__d1, U__d0, P[21]);
  U4DPPG_20_1 U20 (P[23], O_R[22], IN1_R[20], U__d1, U__d0, P[22]);
  U4DPPG_21_1 U21 (P[24], O_R[23], IN1_R[21], U__d1, U__d0, P[23]);
  U4DPPG_22_1 U22 (P[25], O_R[24], IN1_R[22], U__d1, U__d0, P[24]);
  U4DPPG_23_1 U23 (P[26], O_R[25], IN1_R[23], U__d1, U__d0, P[25]);
  U4DPPG_24_1 U24 (P[27], O_R[26], IN1_R[24], U__d1, U__d0, P[26]);
  U4DPPG_25_1 U25 (P[28], O_R[27], IN1_R[25], U__d1, U__d0, P[27]);
  U4DPPG_26_1 U26 (P[29], O_R[28], IN1_R[26], U__d1, U__d0, P[28]);
  U4DPPG_27_1 U27 (P[30], O_R[29], IN1_R[27], U__d1, U__d0, P[29]);
  U4DPPG_28_1 U28 (P[31], O_R[30], IN1_R[28], U__d1, U__d0, P[30]);
  U4DPPG_29_1 U29 (P[32], O_R[31], IN1_R[29], U__d1, U__d0, P[31]);
  U4DPPG_30_1 U30 (P[33], O_R[32], IN1_R[30], U__d1, U__d0, P[32]);
  U4DPPG_31_1 U31 (P[34], O_R[33], IN1_R[31], U__d1, U__d0, P[33]);
  U4DPPG_32_1 U32 (P[35], O_R[34], IN1_R[32], U__d1, U__d0, P[34]);
  U4DPPG_33_1 U33 (P[36], O_R[35], IN1_R[33], U__d1, U__d0, P[35]);
  U4DPPG_34_1 U34 (P[37], O_R[36], IN1_R[34], U__d1, U__d0, P[36]);
  U4DPPG_35_1 U35 (P[38], O_R[37], IN1_R[35], U__d1, U__d0, P[37]);
  U4DPPG_36_1 U36 (P[39], O_R[38], IN1_R[36], U__d1, U__d0, P[38]);
  U4DPPG_37_1 U37 (P[40], O_R[39], IN1_R[37], U__d1, U__d0, P[39]);
  U4DPPG_38_1 U38 (P[41], O_R[40], IN1_R[38], U__d1, U__d0, P[40]);
  U4DPPG_39_1 U39 (P[42], O_R[41], IN1_R[39], U__d1, U__d0, P[41]);
  U4DPPG_40_1 U40 (P[43], O_R[42], IN1_R[40], U__d1, U__d0, P[42]);
  U4DPPG_41_1 U41 (P[44], O_R[43], IN1_R[41], U__d1, U__d0, P[43]);
  U4DPPG_42_1 U42 (P[45], O_R[44], IN1_R[42], U__d1, U__d0, P[44]);
  U4DPPG_43_1 U43 (P[46], O_R[45], IN1_R[43], U__d1, U__d0, P[45]);
  U4DPPG_44_1 U44 (P[47], O_R[46], IN1_R[44], U__d1, U__d0, P[46]);
  U4DPPG_45_1 U45 (P[48], O_R[47], IN1_R[45], U__d1, U__d0, P[47]);
  U4DPPG_46_1 U46 (P[49], O_R[48], IN1_R[46], U__d1, U__d0, P[48]);
  U4DPPG_47_1 U47 (P[50], O_R[49], IN1_R[47], U__d1, U__d0, P[49]);
  U4DPPG_48_1 U48 (P[51], O_R[50], IN1_R[48], U__d1, U__d0, P[50]);
  U4DPPG_49_1 U49 (P[52], O_R[51], IN1_R[49], U__d1, U__d0, P[51]);
  U4DPPG_50_1 U50 (P[53], O_R[52], IN1_R[50], U__d1, U__d0, P[52]);
  U4DPPG_51_1 U51 (P[54], O_R[53], IN1_R[51], U__d1, U__d0, P[53]);
  U4DPPG_52_1 U52 (P[55], O_R[54], IN1_R[52], U__d1, U__d0, P[54]);
  U4DPPG_53_1 U53 (P[56], O_R[55], IN1_R[53], U__d1, U__d0, P[55]);
  U4DPPG_54_1 U54 (P[57], O_R[56], IN1_R[54], U__d1, U__d0, P[56]);
  U4DPPG_55_1 U55 (P[58], O_R[57], IN1_R[55], U__d1, U__d0, P[57]);
  U4DPPG_56_1 U56 (P[59], O_R[58], IN1_R[56], U__d1, U__d0, P[58]);
  U4DPPG_57_1 U57 (P[60], O_R[59], IN1_R[57], U__d1, U__d0, P[59]);
  U4DPPG_58_1 U58 (P[61], O_R[60], IN1_R[58], U__d1, U__d0, P[60]);
  U4DPPG_59_1 U59 (P[62], O_R[61], IN1_R[59], U__d1, U__d0, P[61]);
  U4DPPG_60_1 U60 (P[63], O_R[62], IN1_R[60], U__d1, U__d0, P[62]);
  U4DPPG_61_1 U61 (P[64], O_R[63], IN1_R[61], U__d1, U__d0, P[63]);
  U4DPPG_62_1 U62 (P[65], O_R[64], IN1_R[62], U__d1, U__d0, P[64]);
  U4DPPGH_63_1 U63 (O_T, O_R[65], IN1_T, U__d1, U__d0, P[65]);
endmodule

module TCU4VPPG_63_0_10 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [83:20] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [83:21] P;
  U4DPPGL_0_10 U0 (P[21], O_R[20], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_10 U1 (P[22], O_R[21], IN1_R[1], U__d1, U__d0, P[21]);
  U4DPPG_2_10 U2 (P[23], O_R[22], IN1_R[2], U__d1, U__d0, P[22]);
  U4DPPG_3_10 U3 (P[24], O_R[23], IN1_R[3], U__d1, U__d0, P[23]);
  U4DPPG_4_10 U4 (P[25], O_R[24], IN1_R[4], U__d1, U__d0, P[24]);
  U4DPPG_5_10 U5 (P[26], O_R[25], IN1_R[5], U__d1, U__d0, P[25]);
  U4DPPG_6_10 U6 (P[27], O_R[26], IN1_R[6], U__d1, U__d0, P[26]);
  U4DPPG_7_10 U7 (P[28], O_R[27], IN1_R[7], U__d1, U__d0, P[27]);
  U4DPPG_8_10 U8 (P[29], O_R[28], IN1_R[8], U__d1, U__d0, P[28]);
  U4DPPG_9_10 U9 (P[30], O_R[29], IN1_R[9], U__d1, U__d0, P[29]);
  U4DPPG_10_10 U10 (P[31], O_R[30], IN1_R[10], U__d1, U__d0, P[30]);
  U4DPPG_11_10 U11 (P[32], O_R[31], IN1_R[11], U__d1, U__d0, P[31]);
  U4DPPG_12_10 U12 (P[33], O_R[32], IN1_R[12], U__d1, U__d0, P[32]);
  U4DPPG_13_10 U13 (P[34], O_R[33], IN1_R[13], U__d1, U__d0, P[33]);
  U4DPPG_14_10 U14 (P[35], O_R[34], IN1_R[14], U__d1, U__d0, P[34]);
  U4DPPG_15_10 U15 (P[36], O_R[35], IN1_R[15], U__d1, U__d0, P[35]);
  U4DPPG_16_10 U16 (P[37], O_R[36], IN1_R[16], U__d1, U__d0, P[36]);
  U4DPPG_17_10 U17 (P[38], O_R[37], IN1_R[17], U__d1, U__d0, P[37]);
  U4DPPG_18_10 U18 (P[39], O_R[38], IN1_R[18], U__d1, U__d0, P[38]);
  U4DPPG_19_10 U19 (P[40], O_R[39], IN1_R[19], U__d1, U__d0, P[39]);
  U4DPPG_20_10 U20 (P[41], O_R[40], IN1_R[20], U__d1, U__d0, P[40]);
  U4DPPG_21_10 U21 (P[42], O_R[41], IN1_R[21], U__d1, U__d0, P[41]);
  U4DPPG_22_10 U22 (P[43], O_R[42], IN1_R[22], U__d1, U__d0, P[42]);
  U4DPPG_23_10 U23 (P[44], O_R[43], IN1_R[23], U__d1, U__d0, P[43]);
  U4DPPG_24_10 U24 (P[45], O_R[44], IN1_R[24], U__d1, U__d0, P[44]);
  U4DPPG_25_10 U25 (P[46], O_R[45], IN1_R[25], U__d1, U__d0, P[45]);
  U4DPPG_26_10 U26 (P[47], O_R[46], IN1_R[26], U__d1, U__d0, P[46]);
  U4DPPG_27_10 U27 (P[48], O_R[47], IN1_R[27], U__d1, U__d0, P[47]);
  U4DPPG_28_10 U28 (P[49], O_R[48], IN1_R[28], U__d1, U__d0, P[48]);
  U4DPPG_29_10 U29 (P[50], O_R[49], IN1_R[29], U__d1, U__d0, P[49]);
  U4DPPG_30_10 U30 (P[51], O_R[50], IN1_R[30], U__d1, U__d0, P[50]);
  U4DPPG_31_10 U31 (P[52], O_R[51], IN1_R[31], U__d1, U__d0, P[51]);
  U4DPPG_32_10 U32 (P[53], O_R[52], IN1_R[32], U__d1, U__d0, P[52]);
  U4DPPG_33_10 U33 (P[54], O_R[53], IN1_R[33], U__d1, U__d0, P[53]);
  U4DPPG_34_10 U34 (P[55], O_R[54], IN1_R[34], U__d1, U__d0, P[54]);
  U4DPPG_35_10 U35 (P[56], O_R[55], IN1_R[35], U__d1, U__d0, P[55]);
  U4DPPG_36_10 U36 (P[57], O_R[56], IN1_R[36], U__d1, U__d0, P[56]);
  U4DPPG_37_10 U37 (P[58], O_R[57], IN1_R[37], U__d1, U__d0, P[57]);
  U4DPPG_38_10 U38 (P[59], O_R[58], IN1_R[38], U__d1, U__d0, P[58]);
  U4DPPG_39_10 U39 (P[60], O_R[59], IN1_R[39], U__d1, U__d0, P[59]);
  U4DPPG_40_10 U40 (P[61], O_R[60], IN1_R[40], U__d1, U__d0, P[60]);
  U4DPPG_41_10 U41 (P[62], O_R[61], IN1_R[41], U__d1, U__d0, P[61]);
  U4DPPG_42_10 U42 (P[63], O_R[62], IN1_R[42], U__d1, U__d0, P[62]);
  U4DPPG_43_10 U43 (P[64], O_R[63], IN1_R[43], U__d1, U__d0, P[63]);
  U4DPPG_44_10 U44 (P[65], O_R[64], IN1_R[44], U__d1, U__d0, P[64]);
  U4DPPG_45_10 U45 (P[66], O_R[65], IN1_R[45], U__d1, U__d0, P[65]);
  U4DPPG_46_10 U46 (P[67], O_R[66], IN1_R[46], U__d1, U__d0, P[66]);
  U4DPPG_47_10 U47 (P[68], O_R[67], IN1_R[47], U__d1, U__d0, P[67]);
  U4DPPG_48_10 U48 (P[69], O_R[68], IN1_R[48], U__d1, U__d0, P[68]);
  U4DPPG_49_10 U49 (P[70], O_R[69], IN1_R[49], U__d1, U__d0, P[69]);
  U4DPPG_50_10 U50 (P[71], O_R[70], IN1_R[50], U__d1, U__d0, P[70]);
  U4DPPG_51_10 U51 (P[72], O_R[71], IN1_R[51], U__d1, U__d0, P[71]);
  U4DPPG_52_10 U52 (P[73], O_R[72], IN1_R[52], U__d1, U__d0, P[72]);
  U4DPPG_53_10 U53 (P[74], O_R[73], IN1_R[53], U__d1, U__d0, P[73]);
  U4DPPG_54_10 U54 (P[75], O_R[74], IN1_R[54], U__d1, U__d0, P[74]);
  U4DPPG_55_10 U55 (P[76], O_R[75], IN1_R[55], U__d1, U__d0, P[75]);
  U4DPPG_56_10 U56 (P[77], O_R[76], IN1_R[56], U__d1, U__d0, P[76]);
  U4DPPG_57_10 U57 (P[78], O_R[77], IN1_R[57], U__d1, U__d0, P[77]);
  U4DPPG_58_10 U58 (P[79], O_R[78], IN1_R[58], U__d1, U__d0, P[78]);
  U4DPPG_59_10 U59 (P[80], O_R[79], IN1_R[59], U__d1, U__d0, P[79]);
  U4DPPG_60_10 U60 (P[81], O_R[80], IN1_R[60], U__d1, U__d0, P[80]);
  U4DPPG_61_10 U61 (P[82], O_R[81], IN1_R[61], U__d1, U__d0, P[81]);
  U4DPPG_62_10 U62 (P[83], O_R[82], IN1_R[62], U__d1, U__d0, P[82]);
  U4DPPGH_63_10 U63 (O_T, O_R[83], IN1_T, U__d1, U__d0, P[83]);
endmodule

module TCU4VPPG_63_0_11 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [85:22] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [85:23] P;
  U4DPPGL_0_11 U0 (P[23], O_R[22], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_11 U1 (P[24], O_R[23], IN1_R[1], U__d1, U__d0, P[23]);
  U4DPPG_2_11 U2 (P[25], O_R[24], IN1_R[2], U__d1, U__d0, P[24]);
  U4DPPG_3_11 U3 (P[26], O_R[25], IN1_R[3], U__d1, U__d0, P[25]);
  U4DPPG_4_11 U4 (P[27], O_R[26], IN1_R[4], U__d1, U__d0, P[26]);
  U4DPPG_5_11 U5 (P[28], O_R[27], IN1_R[5], U__d1, U__d0, P[27]);
  U4DPPG_6_11 U6 (P[29], O_R[28], IN1_R[6], U__d1, U__d0, P[28]);
  U4DPPG_7_11 U7 (P[30], O_R[29], IN1_R[7], U__d1, U__d0, P[29]);
  U4DPPG_8_11 U8 (P[31], O_R[30], IN1_R[8], U__d1, U__d0, P[30]);
  U4DPPG_9_11 U9 (P[32], O_R[31], IN1_R[9], U__d1, U__d0, P[31]);
  U4DPPG_10_11 U10 (P[33], O_R[32], IN1_R[10], U__d1, U__d0, P[32]);
  U4DPPG_11_11 U11 (P[34], O_R[33], IN1_R[11], U__d1, U__d0, P[33]);
  U4DPPG_12_11 U12 (P[35], O_R[34], IN1_R[12], U__d1, U__d0, P[34]);
  U4DPPG_13_11 U13 (P[36], O_R[35], IN1_R[13], U__d1, U__d0, P[35]);
  U4DPPG_14_11 U14 (P[37], O_R[36], IN1_R[14], U__d1, U__d0, P[36]);
  U4DPPG_15_11 U15 (P[38], O_R[37], IN1_R[15], U__d1, U__d0, P[37]);
  U4DPPG_16_11 U16 (P[39], O_R[38], IN1_R[16], U__d1, U__d0, P[38]);
  U4DPPG_17_11 U17 (P[40], O_R[39], IN1_R[17], U__d1, U__d0, P[39]);
  U4DPPG_18_11 U18 (P[41], O_R[40], IN1_R[18], U__d1, U__d0, P[40]);
  U4DPPG_19_11 U19 (P[42], O_R[41], IN1_R[19], U__d1, U__d0, P[41]);
  U4DPPG_20_11 U20 (P[43], O_R[42], IN1_R[20], U__d1, U__d0, P[42]);
  U4DPPG_21_11 U21 (P[44], O_R[43], IN1_R[21], U__d1, U__d0, P[43]);
  U4DPPG_22_11 U22 (P[45], O_R[44], IN1_R[22], U__d1, U__d0, P[44]);
  U4DPPG_23_11 U23 (P[46], O_R[45], IN1_R[23], U__d1, U__d0, P[45]);
  U4DPPG_24_11 U24 (P[47], O_R[46], IN1_R[24], U__d1, U__d0, P[46]);
  U4DPPG_25_11 U25 (P[48], O_R[47], IN1_R[25], U__d1, U__d0, P[47]);
  U4DPPG_26_11 U26 (P[49], O_R[48], IN1_R[26], U__d1, U__d0, P[48]);
  U4DPPG_27_11 U27 (P[50], O_R[49], IN1_R[27], U__d1, U__d0, P[49]);
  U4DPPG_28_11 U28 (P[51], O_R[50], IN1_R[28], U__d1, U__d0, P[50]);
  U4DPPG_29_11 U29 (P[52], O_R[51], IN1_R[29], U__d1, U__d0, P[51]);
  U4DPPG_30_11 U30 (P[53], O_R[52], IN1_R[30], U__d1, U__d0, P[52]);
  U4DPPG_31_11 U31 (P[54], O_R[53], IN1_R[31], U__d1, U__d0, P[53]);
  U4DPPG_32_11 U32 (P[55], O_R[54], IN1_R[32], U__d1, U__d0, P[54]);
  U4DPPG_33_11 U33 (P[56], O_R[55], IN1_R[33], U__d1, U__d0, P[55]);
  U4DPPG_34_11 U34 (P[57], O_R[56], IN1_R[34], U__d1, U__d0, P[56]);
  U4DPPG_35_11 U35 (P[58], O_R[57], IN1_R[35], U__d1, U__d0, P[57]);
  U4DPPG_36_11 U36 (P[59], O_R[58], IN1_R[36], U__d1, U__d0, P[58]);
  U4DPPG_37_11 U37 (P[60], O_R[59], IN1_R[37], U__d1, U__d0, P[59]);
  U4DPPG_38_11 U38 (P[61], O_R[60], IN1_R[38], U__d1, U__d0, P[60]);
  U4DPPG_39_11 U39 (P[62], O_R[61], IN1_R[39], U__d1, U__d0, P[61]);
  U4DPPG_40_11 U40 (P[63], O_R[62], IN1_R[40], U__d1, U__d0, P[62]);
  U4DPPG_41_11 U41 (P[64], O_R[63], IN1_R[41], U__d1, U__d0, P[63]);
  U4DPPG_42_11 U42 (P[65], O_R[64], IN1_R[42], U__d1, U__d0, P[64]);
  U4DPPG_43_11 U43 (P[66], O_R[65], IN1_R[43], U__d1, U__d0, P[65]);
  U4DPPG_44_11 U44 (P[67], O_R[66], IN1_R[44], U__d1, U__d0, P[66]);
  U4DPPG_45_11 U45 (P[68], O_R[67], IN1_R[45], U__d1, U__d0, P[67]);
  U4DPPG_46_11 U46 (P[69], O_R[68], IN1_R[46], U__d1, U__d0, P[68]);
  U4DPPG_47_11 U47 (P[70], O_R[69], IN1_R[47], U__d1, U__d0, P[69]);
  U4DPPG_48_11 U48 (P[71], O_R[70], IN1_R[48], U__d1, U__d0, P[70]);
  U4DPPG_49_11 U49 (P[72], O_R[71], IN1_R[49], U__d1, U__d0, P[71]);
  U4DPPG_50_11 U50 (P[73], O_R[72], IN1_R[50], U__d1, U__d0, P[72]);
  U4DPPG_51_11 U51 (P[74], O_R[73], IN1_R[51], U__d1, U__d0, P[73]);
  U4DPPG_52_11 U52 (P[75], O_R[74], IN1_R[52], U__d1, U__d0, P[74]);
  U4DPPG_53_11 U53 (P[76], O_R[75], IN1_R[53], U__d1, U__d0, P[75]);
  U4DPPG_54_11 U54 (P[77], O_R[76], IN1_R[54], U__d1, U__d0, P[76]);
  U4DPPG_55_11 U55 (P[78], O_R[77], IN1_R[55], U__d1, U__d0, P[77]);
  U4DPPG_56_11 U56 (P[79], O_R[78], IN1_R[56], U__d1, U__d0, P[78]);
  U4DPPG_57_11 U57 (P[80], O_R[79], IN1_R[57], U__d1, U__d0, P[79]);
  U4DPPG_58_11 U58 (P[81], O_R[80], IN1_R[58], U__d1, U__d0, P[80]);
  U4DPPG_59_11 U59 (P[82], O_R[81], IN1_R[59], U__d1, U__d0, P[81]);
  U4DPPG_60_11 U60 (P[83], O_R[82], IN1_R[60], U__d1, U__d0, P[82]);
  U4DPPG_61_11 U61 (P[84], O_R[83], IN1_R[61], U__d1, U__d0, P[83]);
  U4DPPG_62_11 U62 (P[85], O_R[84], IN1_R[62], U__d1, U__d0, P[84]);
  U4DPPGH_63_11 U63 (O_T, O_R[85], IN1_T, U__d1, U__d0, P[85]);
endmodule

module TCU4VPPG_63_0_12 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [87:24] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [87:25] P;
  U4DPPGL_0_12 U0 (P[25], O_R[24], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_12 U1 (P[26], O_R[25], IN1_R[1], U__d1, U__d0, P[25]);
  U4DPPG_2_12 U2 (P[27], O_R[26], IN1_R[2], U__d1, U__d0, P[26]);
  U4DPPG_3_12 U3 (P[28], O_R[27], IN1_R[3], U__d1, U__d0, P[27]);
  U4DPPG_4_12 U4 (P[29], O_R[28], IN1_R[4], U__d1, U__d0, P[28]);
  U4DPPG_5_12 U5 (P[30], O_R[29], IN1_R[5], U__d1, U__d0, P[29]);
  U4DPPG_6_12 U6 (P[31], O_R[30], IN1_R[6], U__d1, U__d0, P[30]);
  U4DPPG_7_12 U7 (P[32], O_R[31], IN1_R[7], U__d1, U__d0, P[31]);
  U4DPPG_8_12 U8 (P[33], O_R[32], IN1_R[8], U__d1, U__d0, P[32]);
  U4DPPG_9_12 U9 (P[34], O_R[33], IN1_R[9], U__d1, U__d0, P[33]);
  U4DPPG_10_12 U10 (P[35], O_R[34], IN1_R[10], U__d1, U__d0, P[34]);
  U4DPPG_11_12 U11 (P[36], O_R[35], IN1_R[11], U__d1, U__d0, P[35]);
  U4DPPG_12_12 U12 (P[37], O_R[36], IN1_R[12], U__d1, U__d0, P[36]);
  U4DPPG_13_12 U13 (P[38], O_R[37], IN1_R[13], U__d1, U__d0, P[37]);
  U4DPPG_14_12 U14 (P[39], O_R[38], IN1_R[14], U__d1, U__d0, P[38]);
  U4DPPG_15_12 U15 (P[40], O_R[39], IN1_R[15], U__d1, U__d0, P[39]);
  U4DPPG_16_12 U16 (P[41], O_R[40], IN1_R[16], U__d1, U__d0, P[40]);
  U4DPPG_17_12 U17 (P[42], O_R[41], IN1_R[17], U__d1, U__d0, P[41]);
  U4DPPG_18_12 U18 (P[43], O_R[42], IN1_R[18], U__d1, U__d0, P[42]);
  U4DPPG_19_12 U19 (P[44], O_R[43], IN1_R[19], U__d1, U__d0, P[43]);
  U4DPPG_20_12 U20 (P[45], O_R[44], IN1_R[20], U__d1, U__d0, P[44]);
  U4DPPG_21_12 U21 (P[46], O_R[45], IN1_R[21], U__d1, U__d0, P[45]);
  U4DPPG_22_12 U22 (P[47], O_R[46], IN1_R[22], U__d1, U__d0, P[46]);
  U4DPPG_23_12 U23 (P[48], O_R[47], IN1_R[23], U__d1, U__d0, P[47]);
  U4DPPG_24_12 U24 (P[49], O_R[48], IN1_R[24], U__d1, U__d0, P[48]);
  U4DPPG_25_12 U25 (P[50], O_R[49], IN1_R[25], U__d1, U__d0, P[49]);
  U4DPPG_26_12 U26 (P[51], O_R[50], IN1_R[26], U__d1, U__d0, P[50]);
  U4DPPG_27_12 U27 (P[52], O_R[51], IN1_R[27], U__d1, U__d0, P[51]);
  U4DPPG_28_12 U28 (P[53], O_R[52], IN1_R[28], U__d1, U__d0, P[52]);
  U4DPPG_29_12 U29 (P[54], O_R[53], IN1_R[29], U__d1, U__d0, P[53]);
  U4DPPG_30_12 U30 (P[55], O_R[54], IN1_R[30], U__d1, U__d0, P[54]);
  U4DPPG_31_12 U31 (P[56], O_R[55], IN1_R[31], U__d1, U__d0, P[55]);
  U4DPPG_32_12 U32 (P[57], O_R[56], IN1_R[32], U__d1, U__d0, P[56]);
  U4DPPG_33_12 U33 (P[58], O_R[57], IN1_R[33], U__d1, U__d0, P[57]);
  U4DPPG_34_12 U34 (P[59], O_R[58], IN1_R[34], U__d1, U__d0, P[58]);
  U4DPPG_35_12 U35 (P[60], O_R[59], IN1_R[35], U__d1, U__d0, P[59]);
  U4DPPG_36_12 U36 (P[61], O_R[60], IN1_R[36], U__d1, U__d0, P[60]);
  U4DPPG_37_12 U37 (P[62], O_R[61], IN1_R[37], U__d1, U__d0, P[61]);
  U4DPPG_38_12 U38 (P[63], O_R[62], IN1_R[38], U__d1, U__d0, P[62]);
  U4DPPG_39_12 U39 (P[64], O_R[63], IN1_R[39], U__d1, U__d0, P[63]);
  U4DPPG_40_12 U40 (P[65], O_R[64], IN1_R[40], U__d1, U__d0, P[64]);
  U4DPPG_41_12 U41 (P[66], O_R[65], IN1_R[41], U__d1, U__d0, P[65]);
  U4DPPG_42_12 U42 (P[67], O_R[66], IN1_R[42], U__d1, U__d0, P[66]);
  U4DPPG_43_12 U43 (P[68], O_R[67], IN1_R[43], U__d1, U__d0, P[67]);
  U4DPPG_44_12 U44 (P[69], O_R[68], IN1_R[44], U__d1, U__d0, P[68]);
  U4DPPG_45_12 U45 (P[70], O_R[69], IN1_R[45], U__d1, U__d0, P[69]);
  U4DPPG_46_12 U46 (P[71], O_R[70], IN1_R[46], U__d1, U__d0, P[70]);
  U4DPPG_47_12 U47 (P[72], O_R[71], IN1_R[47], U__d1, U__d0, P[71]);
  U4DPPG_48_12 U48 (P[73], O_R[72], IN1_R[48], U__d1, U__d0, P[72]);
  U4DPPG_49_12 U49 (P[74], O_R[73], IN1_R[49], U__d1, U__d0, P[73]);
  U4DPPG_50_12 U50 (P[75], O_R[74], IN1_R[50], U__d1, U__d0, P[74]);
  U4DPPG_51_12 U51 (P[76], O_R[75], IN1_R[51], U__d1, U__d0, P[75]);
  U4DPPG_52_12 U52 (P[77], O_R[76], IN1_R[52], U__d1, U__d0, P[76]);
  U4DPPG_53_12 U53 (P[78], O_R[77], IN1_R[53], U__d1, U__d0, P[77]);
  U4DPPG_54_12 U54 (P[79], O_R[78], IN1_R[54], U__d1, U__d0, P[78]);
  U4DPPG_55_12 U55 (P[80], O_R[79], IN1_R[55], U__d1, U__d0, P[79]);
  U4DPPG_56_12 U56 (P[81], O_R[80], IN1_R[56], U__d1, U__d0, P[80]);
  U4DPPG_57_12 U57 (P[82], O_R[81], IN1_R[57], U__d1, U__d0, P[81]);
  U4DPPG_58_12 U58 (P[83], O_R[82], IN1_R[58], U__d1, U__d0, P[82]);
  U4DPPG_59_12 U59 (P[84], O_R[83], IN1_R[59], U__d1, U__d0, P[83]);
  U4DPPG_60_12 U60 (P[85], O_R[84], IN1_R[60], U__d1, U__d0, P[84]);
  U4DPPG_61_12 U61 (P[86], O_R[85], IN1_R[61], U__d1, U__d0, P[85]);
  U4DPPG_62_12 U62 (P[87], O_R[86], IN1_R[62], U__d1, U__d0, P[86]);
  U4DPPGH_63_12 U63 (O_T, O_R[87], IN1_T, U__d1, U__d0, P[87]);
endmodule

module TCU4VPPG_63_0_13 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [89:26] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [89:27] P;
  U4DPPGL_0_13 U0 (P[27], O_R[26], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_13 U1 (P[28], O_R[27], IN1_R[1], U__d1, U__d0, P[27]);
  U4DPPG_2_13 U2 (P[29], O_R[28], IN1_R[2], U__d1, U__d0, P[28]);
  U4DPPG_3_13 U3 (P[30], O_R[29], IN1_R[3], U__d1, U__d0, P[29]);
  U4DPPG_4_13 U4 (P[31], O_R[30], IN1_R[4], U__d1, U__d0, P[30]);
  U4DPPG_5_13 U5 (P[32], O_R[31], IN1_R[5], U__d1, U__d0, P[31]);
  U4DPPG_6_13 U6 (P[33], O_R[32], IN1_R[6], U__d1, U__d0, P[32]);
  U4DPPG_7_13 U7 (P[34], O_R[33], IN1_R[7], U__d1, U__d0, P[33]);
  U4DPPG_8_13 U8 (P[35], O_R[34], IN1_R[8], U__d1, U__d0, P[34]);
  U4DPPG_9_13 U9 (P[36], O_R[35], IN1_R[9], U__d1, U__d0, P[35]);
  U4DPPG_10_13 U10 (P[37], O_R[36], IN1_R[10], U__d1, U__d0, P[36]);
  U4DPPG_11_13 U11 (P[38], O_R[37], IN1_R[11], U__d1, U__d0, P[37]);
  U4DPPG_12_13 U12 (P[39], O_R[38], IN1_R[12], U__d1, U__d0, P[38]);
  U4DPPG_13_13 U13 (P[40], O_R[39], IN1_R[13], U__d1, U__d0, P[39]);
  U4DPPG_14_13 U14 (P[41], O_R[40], IN1_R[14], U__d1, U__d0, P[40]);
  U4DPPG_15_13 U15 (P[42], O_R[41], IN1_R[15], U__d1, U__d0, P[41]);
  U4DPPG_16_13 U16 (P[43], O_R[42], IN1_R[16], U__d1, U__d0, P[42]);
  U4DPPG_17_13 U17 (P[44], O_R[43], IN1_R[17], U__d1, U__d0, P[43]);
  U4DPPG_18_13 U18 (P[45], O_R[44], IN1_R[18], U__d1, U__d0, P[44]);
  U4DPPG_19_13 U19 (P[46], O_R[45], IN1_R[19], U__d1, U__d0, P[45]);
  U4DPPG_20_13 U20 (P[47], O_R[46], IN1_R[20], U__d1, U__d0, P[46]);
  U4DPPG_21_13 U21 (P[48], O_R[47], IN1_R[21], U__d1, U__d0, P[47]);
  U4DPPG_22_13 U22 (P[49], O_R[48], IN1_R[22], U__d1, U__d0, P[48]);
  U4DPPG_23_13 U23 (P[50], O_R[49], IN1_R[23], U__d1, U__d0, P[49]);
  U4DPPG_24_13 U24 (P[51], O_R[50], IN1_R[24], U__d1, U__d0, P[50]);
  U4DPPG_25_13 U25 (P[52], O_R[51], IN1_R[25], U__d1, U__d0, P[51]);
  U4DPPG_26_13 U26 (P[53], O_R[52], IN1_R[26], U__d1, U__d0, P[52]);
  U4DPPG_27_13 U27 (P[54], O_R[53], IN1_R[27], U__d1, U__d0, P[53]);
  U4DPPG_28_13 U28 (P[55], O_R[54], IN1_R[28], U__d1, U__d0, P[54]);
  U4DPPG_29_13 U29 (P[56], O_R[55], IN1_R[29], U__d1, U__d0, P[55]);
  U4DPPG_30_13 U30 (P[57], O_R[56], IN1_R[30], U__d1, U__d0, P[56]);
  U4DPPG_31_13 U31 (P[58], O_R[57], IN1_R[31], U__d1, U__d0, P[57]);
  U4DPPG_32_13 U32 (P[59], O_R[58], IN1_R[32], U__d1, U__d0, P[58]);
  U4DPPG_33_13 U33 (P[60], O_R[59], IN1_R[33], U__d1, U__d0, P[59]);
  U4DPPG_34_13 U34 (P[61], O_R[60], IN1_R[34], U__d1, U__d0, P[60]);
  U4DPPG_35_13 U35 (P[62], O_R[61], IN1_R[35], U__d1, U__d0, P[61]);
  U4DPPG_36_13 U36 (P[63], O_R[62], IN1_R[36], U__d1, U__d0, P[62]);
  U4DPPG_37_13 U37 (P[64], O_R[63], IN1_R[37], U__d1, U__d0, P[63]);
  U4DPPG_38_13 U38 (P[65], O_R[64], IN1_R[38], U__d1, U__d0, P[64]);
  U4DPPG_39_13 U39 (P[66], O_R[65], IN1_R[39], U__d1, U__d0, P[65]);
  U4DPPG_40_13 U40 (P[67], O_R[66], IN1_R[40], U__d1, U__d0, P[66]);
  U4DPPG_41_13 U41 (P[68], O_R[67], IN1_R[41], U__d1, U__d0, P[67]);
  U4DPPG_42_13 U42 (P[69], O_R[68], IN1_R[42], U__d1, U__d0, P[68]);
  U4DPPG_43_13 U43 (P[70], O_R[69], IN1_R[43], U__d1, U__d0, P[69]);
  U4DPPG_44_13 U44 (P[71], O_R[70], IN1_R[44], U__d1, U__d0, P[70]);
  U4DPPG_45_13 U45 (P[72], O_R[71], IN1_R[45], U__d1, U__d0, P[71]);
  U4DPPG_46_13 U46 (P[73], O_R[72], IN1_R[46], U__d1, U__d0, P[72]);
  U4DPPG_47_13 U47 (P[74], O_R[73], IN1_R[47], U__d1, U__d0, P[73]);
  U4DPPG_48_13 U48 (P[75], O_R[74], IN1_R[48], U__d1, U__d0, P[74]);
  U4DPPG_49_13 U49 (P[76], O_R[75], IN1_R[49], U__d1, U__d0, P[75]);
  U4DPPG_50_13 U50 (P[77], O_R[76], IN1_R[50], U__d1, U__d0, P[76]);
  U4DPPG_51_13 U51 (P[78], O_R[77], IN1_R[51], U__d1, U__d0, P[77]);
  U4DPPG_52_13 U52 (P[79], O_R[78], IN1_R[52], U__d1, U__d0, P[78]);
  U4DPPG_53_13 U53 (P[80], O_R[79], IN1_R[53], U__d1, U__d0, P[79]);
  U4DPPG_54_13 U54 (P[81], O_R[80], IN1_R[54], U__d1, U__d0, P[80]);
  U4DPPG_55_13 U55 (P[82], O_R[81], IN1_R[55], U__d1, U__d0, P[81]);
  U4DPPG_56_13 U56 (P[83], O_R[82], IN1_R[56], U__d1, U__d0, P[82]);
  U4DPPG_57_13 U57 (P[84], O_R[83], IN1_R[57], U__d1, U__d0, P[83]);
  U4DPPG_58_13 U58 (P[85], O_R[84], IN1_R[58], U__d1, U__d0, P[84]);
  U4DPPG_59_13 U59 (P[86], O_R[85], IN1_R[59], U__d1, U__d0, P[85]);
  U4DPPG_60_13 U60 (P[87], O_R[86], IN1_R[60], U__d1, U__d0, P[86]);
  U4DPPG_61_13 U61 (P[88], O_R[87], IN1_R[61], U__d1, U__d0, P[87]);
  U4DPPG_62_13 U62 (P[89], O_R[88], IN1_R[62], U__d1, U__d0, P[88]);
  U4DPPGH_63_13 U63 (O_T, O_R[89], IN1_T, U__d1, U__d0, P[89]);
endmodule

module TCU4VPPG_63_0_14 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [91:28] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [91:29] P;
  U4DPPGL_0_14 U0 (P[29], O_R[28], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_14 U1 (P[30], O_R[29], IN1_R[1], U__d1, U__d0, P[29]);
  U4DPPG_2_14 U2 (P[31], O_R[30], IN1_R[2], U__d1, U__d0, P[30]);
  U4DPPG_3_14 U3 (P[32], O_R[31], IN1_R[3], U__d1, U__d0, P[31]);
  U4DPPG_4_14 U4 (P[33], O_R[32], IN1_R[4], U__d1, U__d0, P[32]);
  U4DPPG_5_14 U5 (P[34], O_R[33], IN1_R[5], U__d1, U__d0, P[33]);
  U4DPPG_6_14 U6 (P[35], O_R[34], IN1_R[6], U__d1, U__d0, P[34]);
  U4DPPG_7_14 U7 (P[36], O_R[35], IN1_R[7], U__d1, U__d0, P[35]);
  U4DPPG_8_14 U8 (P[37], O_R[36], IN1_R[8], U__d1, U__d0, P[36]);
  U4DPPG_9_14 U9 (P[38], O_R[37], IN1_R[9], U__d1, U__d0, P[37]);
  U4DPPG_10_14 U10 (P[39], O_R[38], IN1_R[10], U__d1, U__d0, P[38]);
  U4DPPG_11_14 U11 (P[40], O_R[39], IN1_R[11], U__d1, U__d0, P[39]);
  U4DPPG_12_14 U12 (P[41], O_R[40], IN1_R[12], U__d1, U__d0, P[40]);
  U4DPPG_13_14 U13 (P[42], O_R[41], IN1_R[13], U__d1, U__d0, P[41]);
  U4DPPG_14_14 U14 (P[43], O_R[42], IN1_R[14], U__d1, U__d0, P[42]);
  U4DPPG_15_14 U15 (P[44], O_R[43], IN1_R[15], U__d1, U__d0, P[43]);
  U4DPPG_16_14 U16 (P[45], O_R[44], IN1_R[16], U__d1, U__d0, P[44]);
  U4DPPG_17_14 U17 (P[46], O_R[45], IN1_R[17], U__d1, U__d0, P[45]);
  U4DPPG_18_14 U18 (P[47], O_R[46], IN1_R[18], U__d1, U__d0, P[46]);
  U4DPPG_19_14 U19 (P[48], O_R[47], IN1_R[19], U__d1, U__d0, P[47]);
  U4DPPG_20_14 U20 (P[49], O_R[48], IN1_R[20], U__d1, U__d0, P[48]);
  U4DPPG_21_14 U21 (P[50], O_R[49], IN1_R[21], U__d1, U__d0, P[49]);
  U4DPPG_22_14 U22 (P[51], O_R[50], IN1_R[22], U__d1, U__d0, P[50]);
  U4DPPG_23_14 U23 (P[52], O_R[51], IN1_R[23], U__d1, U__d0, P[51]);
  U4DPPG_24_14 U24 (P[53], O_R[52], IN1_R[24], U__d1, U__d0, P[52]);
  U4DPPG_25_14 U25 (P[54], O_R[53], IN1_R[25], U__d1, U__d0, P[53]);
  U4DPPG_26_14 U26 (P[55], O_R[54], IN1_R[26], U__d1, U__d0, P[54]);
  U4DPPG_27_14 U27 (P[56], O_R[55], IN1_R[27], U__d1, U__d0, P[55]);
  U4DPPG_28_14 U28 (P[57], O_R[56], IN1_R[28], U__d1, U__d0, P[56]);
  U4DPPG_29_14 U29 (P[58], O_R[57], IN1_R[29], U__d1, U__d0, P[57]);
  U4DPPG_30_14 U30 (P[59], O_R[58], IN1_R[30], U__d1, U__d0, P[58]);
  U4DPPG_31_14 U31 (P[60], O_R[59], IN1_R[31], U__d1, U__d0, P[59]);
  U4DPPG_32_14 U32 (P[61], O_R[60], IN1_R[32], U__d1, U__d0, P[60]);
  U4DPPG_33_14 U33 (P[62], O_R[61], IN1_R[33], U__d1, U__d0, P[61]);
  U4DPPG_34_14 U34 (P[63], O_R[62], IN1_R[34], U__d1, U__d0, P[62]);
  U4DPPG_35_14 U35 (P[64], O_R[63], IN1_R[35], U__d1, U__d0, P[63]);
  U4DPPG_36_14 U36 (P[65], O_R[64], IN1_R[36], U__d1, U__d0, P[64]);
  U4DPPG_37_14 U37 (P[66], O_R[65], IN1_R[37], U__d1, U__d0, P[65]);
  U4DPPG_38_14 U38 (P[67], O_R[66], IN1_R[38], U__d1, U__d0, P[66]);
  U4DPPG_39_14 U39 (P[68], O_R[67], IN1_R[39], U__d1, U__d0, P[67]);
  U4DPPG_40_14 U40 (P[69], O_R[68], IN1_R[40], U__d1, U__d0, P[68]);
  U4DPPG_41_14 U41 (P[70], O_R[69], IN1_R[41], U__d1, U__d0, P[69]);
  U4DPPG_42_14 U42 (P[71], O_R[70], IN1_R[42], U__d1, U__d0, P[70]);
  U4DPPG_43_14 U43 (P[72], O_R[71], IN1_R[43], U__d1, U__d0, P[71]);
  U4DPPG_44_14 U44 (P[73], O_R[72], IN1_R[44], U__d1, U__d0, P[72]);
  U4DPPG_45_14 U45 (P[74], O_R[73], IN1_R[45], U__d1, U__d0, P[73]);
  U4DPPG_46_14 U46 (P[75], O_R[74], IN1_R[46], U__d1, U__d0, P[74]);
  U4DPPG_47_14 U47 (P[76], O_R[75], IN1_R[47], U__d1, U__d0, P[75]);
  U4DPPG_48_14 U48 (P[77], O_R[76], IN1_R[48], U__d1, U__d0, P[76]);
  U4DPPG_49_14 U49 (P[78], O_R[77], IN1_R[49], U__d1, U__d0, P[77]);
  U4DPPG_50_14 U50 (P[79], O_R[78], IN1_R[50], U__d1, U__d0, P[78]);
  U4DPPG_51_14 U51 (P[80], O_R[79], IN1_R[51], U__d1, U__d0, P[79]);
  U4DPPG_52_14 U52 (P[81], O_R[80], IN1_R[52], U__d1, U__d0, P[80]);
  U4DPPG_53_14 U53 (P[82], O_R[81], IN1_R[53], U__d1, U__d0, P[81]);
  U4DPPG_54_14 U54 (P[83], O_R[82], IN1_R[54], U__d1, U__d0, P[82]);
  U4DPPG_55_14 U55 (P[84], O_R[83], IN1_R[55], U__d1, U__d0, P[83]);
  U4DPPG_56_14 U56 (P[85], O_R[84], IN1_R[56], U__d1, U__d0, P[84]);
  U4DPPG_57_14 U57 (P[86], O_R[85], IN1_R[57], U__d1, U__d0, P[85]);
  U4DPPG_58_14 U58 (P[87], O_R[86], IN1_R[58], U__d1, U__d0, P[86]);
  U4DPPG_59_14 U59 (P[88], O_R[87], IN1_R[59], U__d1, U__d0, P[87]);
  U4DPPG_60_14 U60 (P[89], O_R[88], IN1_R[60], U__d1, U__d0, P[88]);
  U4DPPG_61_14 U61 (P[90], O_R[89], IN1_R[61], U__d1, U__d0, P[89]);
  U4DPPG_62_14 U62 (P[91], O_R[90], IN1_R[62], U__d1, U__d0, P[90]);
  U4DPPGH_63_14 U63 (O_T, O_R[91], IN1_T, U__d1, U__d0, P[91]);
endmodule

module TCU4VPPG_63_0_15 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [93:30] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [93:31] P;
  U4DPPGL_0_15 U0 (P[31], O_R[30], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_15 U1 (P[32], O_R[31], IN1_R[1], U__d1, U__d0, P[31]);
  U4DPPG_2_15 U2 (P[33], O_R[32], IN1_R[2], U__d1, U__d0, P[32]);
  U4DPPG_3_15 U3 (P[34], O_R[33], IN1_R[3], U__d1, U__d0, P[33]);
  U4DPPG_4_15 U4 (P[35], O_R[34], IN1_R[4], U__d1, U__d0, P[34]);
  U4DPPG_5_15 U5 (P[36], O_R[35], IN1_R[5], U__d1, U__d0, P[35]);
  U4DPPG_6_15 U6 (P[37], O_R[36], IN1_R[6], U__d1, U__d0, P[36]);
  U4DPPG_7_15 U7 (P[38], O_R[37], IN1_R[7], U__d1, U__d0, P[37]);
  U4DPPG_8_15 U8 (P[39], O_R[38], IN1_R[8], U__d1, U__d0, P[38]);
  U4DPPG_9_15 U9 (P[40], O_R[39], IN1_R[9], U__d1, U__d0, P[39]);
  U4DPPG_10_15 U10 (P[41], O_R[40], IN1_R[10], U__d1, U__d0, P[40]);
  U4DPPG_11_15 U11 (P[42], O_R[41], IN1_R[11], U__d1, U__d0, P[41]);
  U4DPPG_12_15 U12 (P[43], O_R[42], IN1_R[12], U__d1, U__d0, P[42]);
  U4DPPG_13_15 U13 (P[44], O_R[43], IN1_R[13], U__d1, U__d0, P[43]);
  U4DPPG_14_15 U14 (P[45], O_R[44], IN1_R[14], U__d1, U__d0, P[44]);
  U4DPPG_15_15 U15 (P[46], O_R[45], IN1_R[15], U__d1, U__d0, P[45]);
  U4DPPG_16_15 U16 (P[47], O_R[46], IN1_R[16], U__d1, U__d0, P[46]);
  U4DPPG_17_15 U17 (P[48], O_R[47], IN1_R[17], U__d1, U__d0, P[47]);
  U4DPPG_18_15 U18 (P[49], O_R[48], IN1_R[18], U__d1, U__d0, P[48]);
  U4DPPG_19_15 U19 (P[50], O_R[49], IN1_R[19], U__d1, U__d0, P[49]);
  U4DPPG_20_15 U20 (P[51], O_R[50], IN1_R[20], U__d1, U__d0, P[50]);
  U4DPPG_21_15 U21 (P[52], O_R[51], IN1_R[21], U__d1, U__d0, P[51]);
  U4DPPG_22_15 U22 (P[53], O_R[52], IN1_R[22], U__d1, U__d0, P[52]);
  U4DPPG_23_15 U23 (P[54], O_R[53], IN1_R[23], U__d1, U__d0, P[53]);
  U4DPPG_24_15 U24 (P[55], O_R[54], IN1_R[24], U__d1, U__d0, P[54]);
  U4DPPG_25_15 U25 (P[56], O_R[55], IN1_R[25], U__d1, U__d0, P[55]);
  U4DPPG_26_15 U26 (P[57], O_R[56], IN1_R[26], U__d1, U__d0, P[56]);
  U4DPPG_27_15 U27 (P[58], O_R[57], IN1_R[27], U__d1, U__d0, P[57]);
  U4DPPG_28_15 U28 (P[59], O_R[58], IN1_R[28], U__d1, U__d0, P[58]);
  U4DPPG_29_15 U29 (P[60], O_R[59], IN1_R[29], U__d1, U__d0, P[59]);
  U4DPPG_30_15 U30 (P[61], O_R[60], IN1_R[30], U__d1, U__d0, P[60]);
  U4DPPG_31_15 U31 (P[62], O_R[61], IN1_R[31], U__d1, U__d0, P[61]);
  U4DPPG_32_15 U32 (P[63], O_R[62], IN1_R[32], U__d1, U__d0, P[62]);
  U4DPPG_33_15 U33 (P[64], O_R[63], IN1_R[33], U__d1, U__d0, P[63]);
  U4DPPG_34_15 U34 (P[65], O_R[64], IN1_R[34], U__d1, U__d0, P[64]);
  U4DPPG_35_15 U35 (P[66], O_R[65], IN1_R[35], U__d1, U__d0, P[65]);
  U4DPPG_36_15 U36 (P[67], O_R[66], IN1_R[36], U__d1, U__d0, P[66]);
  U4DPPG_37_15 U37 (P[68], O_R[67], IN1_R[37], U__d1, U__d0, P[67]);
  U4DPPG_38_15 U38 (P[69], O_R[68], IN1_R[38], U__d1, U__d0, P[68]);
  U4DPPG_39_15 U39 (P[70], O_R[69], IN1_R[39], U__d1, U__d0, P[69]);
  U4DPPG_40_15 U40 (P[71], O_R[70], IN1_R[40], U__d1, U__d0, P[70]);
  U4DPPG_41_15 U41 (P[72], O_R[71], IN1_R[41], U__d1, U__d0, P[71]);
  U4DPPG_42_15 U42 (P[73], O_R[72], IN1_R[42], U__d1, U__d0, P[72]);
  U4DPPG_43_15 U43 (P[74], O_R[73], IN1_R[43], U__d1, U__d0, P[73]);
  U4DPPG_44_15 U44 (P[75], O_R[74], IN1_R[44], U__d1, U__d0, P[74]);
  U4DPPG_45_15 U45 (P[76], O_R[75], IN1_R[45], U__d1, U__d0, P[75]);
  U4DPPG_46_15 U46 (P[77], O_R[76], IN1_R[46], U__d1, U__d0, P[76]);
  U4DPPG_47_15 U47 (P[78], O_R[77], IN1_R[47], U__d1, U__d0, P[77]);
  U4DPPG_48_15 U48 (P[79], O_R[78], IN1_R[48], U__d1, U__d0, P[78]);
  U4DPPG_49_15 U49 (P[80], O_R[79], IN1_R[49], U__d1, U__d0, P[79]);
  U4DPPG_50_15 U50 (P[81], O_R[80], IN1_R[50], U__d1, U__d0, P[80]);
  U4DPPG_51_15 U51 (P[82], O_R[81], IN1_R[51], U__d1, U__d0, P[81]);
  U4DPPG_52_15 U52 (P[83], O_R[82], IN1_R[52], U__d1, U__d0, P[82]);
  U4DPPG_53_15 U53 (P[84], O_R[83], IN1_R[53], U__d1, U__d0, P[83]);
  U4DPPG_54_15 U54 (P[85], O_R[84], IN1_R[54], U__d1, U__d0, P[84]);
  U4DPPG_55_15 U55 (P[86], O_R[85], IN1_R[55], U__d1, U__d0, P[85]);
  U4DPPG_56_15 U56 (P[87], O_R[86], IN1_R[56], U__d1, U__d0, P[86]);
  U4DPPG_57_15 U57 (P[88], O_R[87], IN1_R[57], U__d1, U__d0, P[87]);
  U4DPPG_58_15 U58 (P[89], O_R[88], IN1_R[58], U__d1, U__d0, P[88]);
  U4DPPG_59_15 U59 (P[90], O_R[89], IN1_R[59], U__d1, U__d0, P[89]);
  U4DPPG_60_15 U60 (P[91], O_R[90], IN1_R[60], U__d1, U__d0, P[90]);
  U4DPPG_61_15 U61 (P[92], O_R[91], IN1_R[61], U__d1, U__d0, P[91]);
  U4DPPG_62_15 U62 (P[93], O_R[92], IN1_R[62], U__d1, U__d0, P[92]);
  U4DPPGH_63_15 U63 (O_T, O_R[93], IN1_T, U__d1, U__d0, P[93]);
endmodule

module TCU4VPPG_63_0_16 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [95:32] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [95:33] P;
  U4DPPGL_0_16 U0 (P[33], O_R[32], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_16 U1 (P[34], O_R[33], IN1_R[1], U__d1, U__d0, P[33]);
  U4DPPG_2_16 U2 (P[35], O_R[34], IN1_R[2], U__d1, U__d0, P[34]);
  U4DPPG_3_16 U3 (P[36], O_R[35], IN1_R[3], U__d1, U__d0, P[35]);
  U4DPPG_4_16 U4 (P[37], O_R[36], IN1_R[4], U__d1, U__d0, P[36]);
  U4DPPG_5_16 U5 (P[38], O_R[37], IN1_R[5], U__d1, U__d0, P[37]);
  U4DPPG_6_16 U6 (P[39], O_R[38], IN1_R[6], U__d1, U__d0, P[38]);
  U4DPPG_7_16 U7 (P[40], O_R[39], IN1_R[7], U__d1, U__d0, P[39]);
  U4DPPG_8_16 U8 (P[41], O_R[40], IN1_R[8], U__d1, U__d0, P[40]);
  U4DPPG_9_16 U9 (P[42], O_R[41], IN1_R[9], U__d1, U__d0, P[41]);
  U4DPPG_10_16 U10 (P[43], O_R[42], IN1_R[10], U__d1, U__d0, P[42]);
  U4DPPG_11_16 U11 (P[44], O_R[43], IN1_R[11], U__d1, U__d0, P[43]);
  U4DPPG_12_16 U12 (P[45], O_R[44], IN1_R[12], U__d1, U__d0, P[44]);
  U4DPPG_13_16 U13 (P[46], O_R[45], IN1_R[13], U__d1, U__d0, P[45]);
  U4DPPG_14_16 U14 (P[47], O_R[46], IN1_R[14], U__d1, U__d0, P[46]);
  U4DPPG_15_16 U15 (P[48], O_R[47], IN1_R[15], U__d1, U__d0, P[47]);
  U4DPPG_16_16 U16 (P[49], O_R[48], IN1_R[16], U__d1, U__d0, P[48]);
  U4DPPG_17_16 U17 (P[50], O_R[49], IN1_R[17], U__d1, U__d0, P[49]);
  U4DPPG_18_16 U18 (P[51], O_R[50], IN1_R[18], U__d1, U__d0, P[50]);
  U4DPPG_19_16 U19 (P[52], O_R[51], IN1_R[19], U__d1, U__d0, P[51]);
  U4DPPG_20_16 U20 (P[53], O_R[52], IN1_R[20], U__d1, U__d0, P[52]);
  U4DPPG_21_16 U21 (P[54], O_R[53], IN1_R[21], U__d1, U__d0, P[53]);
  U4DPPG_22_16 U22 (P[55], O_R[54], IN1_R[22], U__d1, U__d0, P[54]);
  U4DPPG_23_16 U23 (P[56], O_R[55], IN1_R[23], U__d1, U__d0, P[55]);
  U4DPPG_24_16 U24 (P[57], O_R[56], IN1_R[24], U__d1, U__d0, P[56]);
  U4DPPG_25_16 U25 (P[58], O_R[57], IN1_R[25], U__d1, U__d0, P[57]);
  U4DPPG_26_16 U26 (P[59], O_R[58], IN1_R[26], U__d1, U__d0, P[58]);
  U4DPPG_27_16 U27 (P[60], O_R[59], IN1_R[27], U__d1, U__d0, P[59]);
  U4DPPG_28_16 U28 (P[61], O_R[60], IN1_R[28], U__d1, U__d0, P[60]);
  U4DPPG_29_16 U29 (P[62], O_R[61], IN1_R[29], U__d1, U__d0, P[61]);
  U4DPPG_30_16 U30 (P[63], O_R[62], IN1_R[30], U__d1, U__d0, P[62]);
  U4DPPG_31_16 U31 (P[64], O_R[63], IN1_R[31], U__d1, U__d0, P[63]);
  U4DPPG_32_16 U32 (P[65], O_R[64], IN1_R[32], U__d1, U__d0, P[64]);
  U4DPPG_33_16 U33 (P[66], O_R[65], IN1_R[33], U__d1, U__d0, P[65]);
  U4DPPG_34_16 U34 (P[67], O_R[66], IN1_R[34], U__d1, U__d0, P[66]);
  U4DPPG_35_16 U35 (P[68], O_R[67], IN1_R[35], U__d1, U__d0, P[67]);
  U4DPPG_36_16 U36 (P[69], O_R[68], IN1_R[36], U__d1, U__d0, P[68]);
  U4DPPG_37_16 U37 (P[70], O_R[69], IN1_R[37], U__d1, U__d0, P[69]);
  U4DPPG_38_16 U38 (P[71], O_R[70], IN1_R[38], U__d1, U__d0, P[70]);
  U4DPPG_39_16 U39 (P[72], O_R[71], IN1_R[39], U__d1, U__d0, P[71]);
  U4DPPG_40_16 U40 (P[73], O_R[72], IN1_R[40], U__d1, U__d0, P[72]);
  U4DPPG_41_16 U41 (P[74], O_R[73], IN1_R[41], U__d1, U__d0, P[73]);
  U4DPPG_42_16 U42 (P[75], O_R[74], IN1_R[42], U__d1, U__d0, P[74]);
  U4DPPG_43_16 U43 (P[76], O_R[75], IN1_R[43], U__d1, U__d0, P[75]);
  U4DPPG_44_16 U44 (P[77], O_R[76], IN1_R[44], U__d1, U__d0, P[76]);
  U4DPPG_45_16 U45 (P[78], O_R[77], IN1_R[45], U__d1, U__d0, P[77]);
  U4DPPG_46_16 U46 (P[79], O_R[78], IN1_R[46], U__d1, U__d0, P[78]);
  U4DPPG_47_16 U47 (P[80], O_R[79], IN1_R[47], U__d1, U__d0, P[79]);
  U4DPPG_48_16 U48 (P[81], O_R[80], IN1_R[48], U__d1, U__d0, P[80]);
  U4DPPG_49_16 U49 (P[82], O_R[81], IN1_R[49], U__d1, U__d0, P[81]);
  U4DPPG_50_16 U50 (P[83], O_R[82], IN1_R[50], U__d1, U__d0, P[82]);
  U4DPPG_51_16 U51 (P[84], O_R[83], IN1_R[51], U__d1, U__d0, P[83]);
  U4DPPG_52_16 U52 (P[85], O_R[84], IN1_R[52], U__d1, U__d0, P[84]);
  U4DPPG_53_16 U53 (P[86], O_R[85], IN1_R[53], U__d1, U__d0, P[85]);
  U4DPPG_54_16 U54 (P[87], O_R[86], IN1_R[54], U__d1, U__d0, P[86]);
  U4DPPG_55_16 U55 (P[88], O_R[87], IN1_R[55], U__d1, U__d0, P[87]);
  U4DPPG_56_16 U56 (P[89], O_R[88], IN1_R[56], U__d1, U__d0, P[88]);
  U4DPPG_57_16 U57 (P[90], O_R[89], IN1_R[57], U__d1, U__d0, P[89]);
  U4DPPG_58_16 U58 (P[91], O_R[90], IN1_R[58], U__d1, U__d0, P[90]);
  U4DPPG_59_16 U59 (P[92], O_R[91], IN1_R[59], U__d1, U__d0, P[91]);
  U4DPPG_60_16 U60 (P[93], O_R[92], IN1_R[60], U__d1, U__d0, P[92]);
  U4DPPG_61_16 U61 (P[94], O_R[93], IN1_R[61], U__d1, U__d0, P[93]);
  U4DPPG_62_16 U62 (P[95], O_R[94], IN1_R[62], U__d1, U__d0, P[94]);
  U4DPPGH_63_16 U63 (O_T, O_R[95], IN1_T, U__d1, U__d0, P[95]);
endmodule

module TCU4VPPG_63_0_17 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [97:34] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [97:35] P;
  U4DPPGL_0_17 U0 (P[35], O_R[34], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_17 U1 (P[36], O_R[35], IN1_R[1], U__d1, U__d0, P[35]);
  U4DPPG_2_17 U2 (P[37], O_R[36], IN1_R[2], U__d1, U__d0, P[36]);
  U4DPPG_3_17 U3 (P[38], O_R[37], IN1_R[3], U__d1, U__d0, P[37]);
  U4DPPG_4_17 U4 (P[39], O_R[38], IN1_R[4], U__d1, U__d0, P[38]);
  U4DPPG_5_17 U5 (P[40], O_R[39], IN1_R[5], U__d1, U__d0, P[39]);
  U4DPPG_6_17 U6 (P[41], O_R[40], IN1_R[6], U__d1, U__d0, P[40]);
  U4DPPG_7_17 U7 (P[42], O_R[41], IN1_R[7], U__d1, U__d0, P[41]);
  U4DPPG_8_17 U8 (P[43], O_R[42], IN1_R[8], U__d1, U__d0, P[42]);
  U4DPPG_9_17 U9 (P[44], O_R[43], IN1_R[9], U__d1, U__d0, P[43]);
  U4DPPG_10_17 U10 (P[45], O_R[44], IN1_R[10], U__d1, U__d0, P[44]);
  U4DPPG_11_17 U11 (P[46], O_R[45], IN1_R[11], U__d1, U__d0, P[45]);
  U4DPPG_12_17 U12 (P[47], O_R[46], IN1_R[12], U__d1, U__d0, P[46]);
  U4DPPG_13_17 U13 (P[48], O_R[47], IN1_R[13], U__d1, U__d0, P[47]);
  U4DPPG_14_17 U14 (P[49], O_R[48], IN1_R[14], U__d1, U__d0, P[48]);
  U4DPPG_15_17 U15 (P[50], O_R[49], IN1_R[15], U__d1, U__d0, P[49]);
  U4DPPG_16_17 U16 (P[51], O_R[50], IN1_R[16], U__d1, U__d0, P[50]);
  U4DPPG_17_17 U17 (P[52], O_R[51], IN1_R[17], U__d1, U__d0, P[51]);
  U4DPPG_18_17 U18 (P[53], O_R[52], IN1_R[18], U__d1, U__d0, P[52]);
  U4DPPG_19_17 U19 (P[54], O_R[53], IN1_R[19], U__d1, U__d0, P[53]);
  U4DPPG_20_17 U20 (P[55], O_R[54], IN1_R[20], U__d1, U__d0, P[54]);
  U4DPPG_21_17 U21 (P[56], O_R[55], IN1_R[21], U__d1, U__d0, P[55]);
  U4DPPG_22_17 U22 (P[57], O_R[56], IN1_R[22], U__d1, U__d0, P[56]);
  U4DPPG_23_17 U23 (P[58], O_R[57], IN1_R[23], U__d1, U__d0, P[57]);
  U4DPPG_24_17 U24 (P[59], O_R[58], IN1_R[24], U__d1, U__d0, P[58]);
  U4DPPG_25_17 U25 (P[60], O_R[59], IN1_R[25], U__d1, U__d0, P[59]);
  U4DPPG_26_17 U26 (P[61], O_R[60], IN1_R[26], U__d1, U__d0, P[60]);
  U4DPPG_27_17 U27 (P[62], O_R[61], IN1_R[27], U__d1, U__d0, P[61]);
  U4DPPG_28_17 U28 (P[63], O_R[62], IN1_R[28], U__d1, U__d0, P[62]);
  U4DPPG_29_17 U29 (P[64], O_R[63], IN1_R[29], U__d1, U__d0, P[63]);
  U4DPPG_30_17 U30 (P[65], O_R[64], IN1_R[30], U__d1, U__d0, P[64]);
  U4DPPG_31_17 U31 (P[66], O_R[65], IN1_R[31], U__d1, U__d0, P[65]);
  U4DPPG_32_17 U32 (P[67], O_R[66], IN1_R[32], U__d1, U__d0, P[66]);
  U4DPPG_33_17 U33 (P[68], O_R[67], IN1_R[33], U__d1, U__d0, P[67]);
  U4DPPG_34_17 U34 (P[69], O_R[68], IN1_R[34], U__d1, U__d0, P[68]);
  U4DPPG_35_17 U35 (P[70], O_R[69], IN1_R[35], U__d1, U__d0, P[69]);
  U4DPPG_36_17 U36 (P[71], O_R[70], IN1_R[36], U__d1, U__d0, P[70]);
  U4DPPG_37_17 U37 (P[72], O_R[71], IN1_R[37], U__d1, U__d0, P[71]);
  U4DPPG_38_17 U38 (P[73], O_R[72], IN1_R[38], U__d1, U__d0, P[72]);
  U4DPPG_39_17 U39 (P[74], O_R[73], IN1_R[39], U__d1, U__d0, P[73]);
  U4DPPG_40_17 U40 (P[75], O_R[74], IN1_R[40], U__d1, U__d0, P[74]);
  U4DPPG_41_17 U41 (P[76], O_R[75], IN1_R[41], U__d1, U__d0, P[75]);
  U4DPPG_42_17 U42 (P[77], O_R[76], IN1_R[42], U__d1, U__d0, P[76]);
  U4DPPG_43_17 U43 (P[78], O_R[77], IN1_R[43], U__d1, U__d0, P[77]);
  U4DPPG_44_17 U44 (P[79], O_R[78], IN1_R[44], U__d1, U__d0, P[78]);
  U4DPPG_45_17 U45 (P[80], O_R[79], IN1_R[45], U__d1, U__d0, P[79]);
  U4DPPG_46_17 U46 (P[81], O_R[80], IN1_R[46], U__d1, U__d0, P[80]);
  U4DPPG_47_17 U47 (P[82], O_R[81], IN1_R[47], U__d1, U__d0, P[81]);
  U4DPPG_48_17 U48 (P[83], O_R[82], IN1_R[48], U__d1, U__d0, P[82]);
  U4DPPG_49_17 U49 (P[84], O_R[83], IN1_R[49], U__d1, U__d0, P[83]);
  U4DPPG_50_17 U50 (P[85], O_R[84], IN1_R[50], U__d1, U__d0, P[84]);
  U4DPPG_51_17 U51 (P[86], O_R[85], IN1_R[51], U__d1, U__d0, P[85]);
  U4DPPG_52_17 U52 (P[87], O_R[86], IN1_R[52], U__d1, U__d0, P[86]);
  U4DPPG_53_17 U53 (P[88], O_R[87], IN1_R[53], U__d1, U__d0, P[87]);
  U4DPPG_54_17 U54 (P[89], O_R[88], IN1_R[54], U__d1, U__d0, P[88]);
  U4DPPG_55_17 U55 (P[90], O_R[89], IN1_R[55], U__d1, U__d0, P[89]);
  U4DPPG_56_17 U56 (P[91], O_R[90], IN1_R[56], U__d1, U__d0, P[90]);
  U4DPPG_57_17 U57 (P[92], O_R[91], IN1_R[57], U__d1, U__d0, P[91]);
  U4DPPG_58_17 U58 (P[93], O_R[92], IN1_R[58], U__d1, U__d0, P[92]);
  U4DPPG_59_17 U59 (P[94], O_R[93], IN1_R[59], U__d1, U__d0, P[93]);
  U4DPPG_60_17 U60 (P[95], O_R[94], IN1_R[60], U__d1, U__d0, P[94]);
  U4DPPG_61_17 U61 (P[96], O_R[95], IN1_R[61], U__d1, U__d0, P[95]);
  U4DPPG_62_17 U62 (P[97], O_R[96], IN1_R[62], U__d1, U__d0, P[96]);
  U4DPPGH_63_17 U63 (O_T, O_R[97], IN1_T, U__d1, U__d0, P[97]);
endmodule

module TCU4VPPG_63_0_18 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [99:36] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [99:37] P;
  U4DPPGL_0_18 U0 (P[37], O_R[36], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_18 U1 (P[38], O_R[37], IN1_R[1], U__d1, U__d0, P[37]);
  U4DPPG_2_18 U2 (P[39], O_R[38], IN1_R[2], U__d1, U__d0, P[38]);
  U4DPPG_3_18 U3 (P[40], O_R[39], IN1_R[3], U__d1, U__d0, P[39]);
  U4DPPG_4_18 U4 (P[41], O_R[40], IN1_R[4], U__d1, U__d0, P[40]);
  U4DPPG_5_18 U5 (P[42], O_R[41], IN1_R[5], U__d1, U__d0, P[41]);
  U4DPPG_6_18 U6 (P[43], O_R[42], IN1_R[6], U__d1, U__d0, P[42]);
  U4DPPG_7_18 U7 (P[44], O_R[43], IN1_R[7], U__d1, U__d0, P[43]);
  U4DPPG_8_18 U8 (P[45], O_R[44], IN1_R[8], U__d1, U__d0, P[44]);
  U4DPPG_9_18 U9 (P[46], O_R[45], IN1_R[9], U__d1, U__d0, P[45]);
  U4DPPG_10_18 U10 (P[47], O_R[46], IN1_R[10], U__d1, U__d0, P[46]);
  U4DPPG_11_18 U11 (P[48], O_R[47], IN1_R[11], U__d1, U__d0, P[47]);
  U4DPPG_12_18 U12 (P[49], O_R[48], IN1_R[12], U__d1, U__d0, P[48]);
  U4DPPG_13_18 U13 (P[50], O_R[49], IN1_R[13], U__d1, U__d0, P[49]);
  U4DPPG_14_18 U14 (P[51], O_R[50], IN1_R[14], U__d1, U__d0, P[50]);
  U4DPPG_15_18 U15 (P[52], O_R[51], IN1_R[15], U__d1, U__d0, P[51]);
  U4DPPG_16_18 U16 (P[53], O_R[52], IN1_R[16], U__d1, U__d0, P[52]);
  U4DPPG_17_18 U17 (P[54], O_R[53], IN1_R[17], U__d1, U__d0, P[53]);
  U4DPPG_18_18 U18 (P[55], O_R[54], IN1_R[18], U__d1, U__d0, P[54]);
  U4DPPG_19_18 U19 (P[56], O_R[55], IN1_R[19], U__d1, U__d0, P[55]);
  U4DPPG_20_18 U20 (P[57], O_R[56], IN1_R[20], U__d1, U__d0, P[56]);
  U4DPPG_21_18 U21 (P[58], O_R[57], IN1_R[21], U__d1, U__d0, P[57]);
  U4DPPG_22_18 U22 (P[59], O_R[58], IN1_R[22], U__d1, U__d0, P[58]);
  U4DPPG_23_18 U23 (P[60], O_R[59], IN1_R[23], U__d1, U__d0, P[59]);
  U4DPPG_24_18 U24 (P[61], O_R[60], IN1_R[24], U__d1, U__d0, P[60]);
  U4DPPG_25_18 U25 (P[62], O_R[61], IN1_R[25], U__d1, U__d0, P[61]);
  U4DPPG_26_18 U26 (P[63], O_R[62], IN1_R[26], U__d1, U__d0, P[62]);
  U4DPPG_27_18 U27 (P[64], O_R[63], IN1_R[27], U__d1, U__d0, P[63]);
  U4DPPG_28_18 U28 (P[65], O_R[64], IN1_R[28], U__d1, U__d0, P[64]);
  U4DPPG_29_18 U29 (P[66], O_R[65], IN1_R[29], U__d1, U__d0, P[65]);
  U4DPPG_30_18 U30 (P[67], O_R[66], IN1_R[30], U__d1, U__d0, P[66]);
  U4DPPG_31_18 U31 (P[68], O_R[67], IN1_R[31], U__d1, U__d0, P[67]);
  U4DPPG_32_18 U32 (P[69], O_R[68], IN1_R[32], U__d1, U__d0, P[68]);
  U4DPPG_33_18 U33 (P[70], O_R[69], IN1_R[33], U__d1, U__d0, P[69]);
  U4DPPG_34_18 U34 (P[71], O_R[70], IN1_R[34], U__d1, U__d0, P[70]);
  U4DPPG_35_18 U35 (P[72], O_R[71], IN1_R[35], U__d1, U__d0, P[71]);
  U4DPPG_36_18 U36 (P[73], O_R[72], IN1_R[36], U__d1, U__d0, P[72]);
  U4DPPG_37_18 U37 (P[74], O_R[73], IN1_R[37], U__d1, U__d0, P[73]);
  U4DPPG_38_18 U38 (P[75], O_R[74], IN1_R[38], U__d1, U__d0, P[74]);
  U4DPPG_39_18 U39 (P[76], O_R[75], IN1_R[39], U__d1, U__d0, P[75]);
  U4DPPG_40_18 U40 (P[77], O_R[76], IN1_R[40], U__d1, U__d0, P[76]);
  U4DPPG_41_18 U41 (P[78], O_R[77], IN1_R[41], U__d1, U__d0, P[77]);
  U4DPPG_42_18 U42 (P[79], O_R[78], IN1_R[42], U__d1, U__d0, P[78]);
  U4DPPG_43_18 U43 (P[80], O_R[79], IN1_R[43], U__d1, U__d0, P[79]);
  U4DPPG_44_18 U44 (P[81], O_R[80], IN1_R[44], U__d1, U__d0, P[80]);
  U4DPPG_45_18 U45 (P[82], O_R[81], IN1_R[45], U__d1, U__d0, P[81]);
  U4DPPG_46_18 U46 (P[83], O_R[82], IN1_R[46], U__d1, U__d0, P[82]);
  U4DPPG_47_18 U47 (P[84], O_R[83], IN1_R[47], U__d1, U__d0, P[83]);
  U4DPPG_48_18 U48 (P[85], O_R[84], IN1_R[48], U__d1, U__d0, P[84]);
  U4DPPG_49_18 U49 (P[86], O_R[85], IN1_R[49], U__d1, U__d0, P[85]);
  U4DPPG_50_18 U50 (P[87], O_R[86], IN1_R[50], U__d1, U__d0, P[86]);
  U4DPPG_51_18 U51 (P[88], O_R[87], IN1_R[51], U__d1, U__d0, P[87]);
  U4DPPG_52_18 U52 (P[89], O_R[88], IN1_R[52], U__d1, U__d0, P[88]);
  U4DPPG_53_18 U53 (P[90], O_R[89], IN1_R[53], U__d1, U__d0, P[89]);
  U4DPPG_54_18 U54 (P[91], O_R[90], IN1_R[54], U__d1, U__d0, P[90]);
  U4DPPG_55_18 U55 (P[92], O_R[91], IN1_R[55], U__d1, U__d0, P[91]);
  U4DPPG_56_18 U56 (P[93], O_R[92], IN1_R[56], U__d1, U__d0, P[92]);
  U4DPPG_57_18 U57 (P[94], O_R[93], IN1_R[57], U__d1, U__d0, P[93]);
  U4DPPG_58_18 U58 (P[95], O_R[94], IN1_R[58], U__d1, U__d0, P[94]);
  U4DPPG_59_18 U59 (P[96], O_R[95], IN1_R[59], U__d1, U__d0, P[95]);
  U4DPPG_60_18 U60 (P[97], O_R[96], IN1_R[60], U__d1, U__d0, P[96]);
  U4DPPG_61_18 U61 (P[98], O_R[97], IN1_R[61], U__d1, U__d0, P[97]);
  U4DPPG_62_18 U62 (P[99], O_R[98], IN1_R[62], U__d1, U__d0, P[98]);
  U4DPPGH_63_18 U63 (O_T, O_R[99], IN1_T, U__d1, U__d0, P[99]);
endmodule

module TCU4VPPG_63_0_19 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [101:38] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [101:39] P;
  U4DPPGL_0_19 U0 (P[39], O_R[38], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_19 U1 (P[40], O_R[39], IN1_R[1], U__d1, U__d0, P[39]);
  U4DPPG_2_19 U2 (P[41], O_R[40], IN1_R[2], U__d1, U__d0, P[40]);
  U4DPPG_3_19 U3 (P[42], O_R[41], IN1_R[3], U__d1, U__d0, P[41]);
  U4DPPG_4_19 U4 (P[43], O_R[42], IN1_R[4], U__d1, U__d0, P[42]);
  U4DPPG_5_19 U5 (P[44], O_R[43], IN1_R[5], U__d1, U__d0, P[43]);
  U4DPPG_6_19 U6 (P[45], O_R[44], IN1_R[6], U__d1, U__d0, P[44]);
  U4DPPG_7_19 U7 (P[46], O_R[45], IN1_R[7], U__d1, U__d0, P[45]);
  U4DPPG_8_19 U8 (P[47], O_R[46], IN1_R[8], U__d1, U__d0, P[46]);
  U4DPPG_9_19 U9 (P[48], O_R[47], IN1_R[9], U__d1, U__d0, P[47]);
  U4DPPG_10_19 U10 (P[49], O_R[48], IN1_R[10], U__d1, U__d0, P[48]);
  U4DPPG_11_19 U11 (P[50], O_R[49], IN1_R[11], U__d1, U__d0, P[49]);
  U4DPPG_12_19 U12 (P[51], O_R[50], IN1_R[12], U__d1, U__d0, P[50]);
  U4DPPG_13_19 U13 (P[52], O_R[51], IN1_R[13], U__d1, U__d0, P[51]);
  U4DPPG_14_19 U14 (P[53], O_R[52], IN1_R[14], U__d1, U__d0, P[52]);
  U4DPPG_15_19 U15 (P[54], O_R[53], IN1_R[15], U__d1, U__d0, P[53]);
  U4DPPG_16_19 U16 (P[55], O_R[54], IN1_R[16], U__d1, U__d0, P[54]);
  U4DPPG_17_19 U17 (P[56], O_R[55], IN1_R[17], U__d1, U__d0, P[55]);
  U4DPPG_18_19 U18 (P[57], O_R[56], IN1_R[18], U__d1, U__d0, P[56]);
  U4DPPG_19_19 U19 (P[58], O_R[57], IN1_R[19], U__d1, U__d0, P[57]);
  U4DPPG_20_19 U20 (P[59], O_R[58], IN1_R[20], U__d1, U__d0, P[58]);
  U4DPPG_21_19 U21 (P[60], O_R[59], IN1_R[21], U__d1, U__d0, P[59]);
  U4DPPG_22_19 U22 (P[61], O_R[60], IN1_R[22], U__d1, U__d0, P[60]);
  U4DPPG_23_19 U23 (P[62], O_R[61], IN1_R[23], U__d1, U__d0, P[61]);
  U4DPPG_24_19 U24 (P[63], O_R[62], IN1_R[24], U__d1, U__d0, P[62]);
  U4DPPG_25_19 U25 (P[64], O_R[63], IN1_R[25], U__d1, U__d0, P[63]);
  U4DPPG_26_19 U26 (P[65], O_R[64], IN1_R[26], U__d1, U__d0, P[64]);
  U4DPPG_27_19 U27 (P[66], O_R[65], IN1_R[27], U__d1, U__d0, P[65]);
  U4DPPG_28_19 U28 (P[67], O_R[66], IN1_R[28], U__d1, U__d0, P[66]);
  U4DPPG_29_19 U29 (P[68], O_R[67], IN1_R[29], U__d1, U__d0, P[67]);
  U4DPPG_30_19 U30 (P[69], O_R[68], IN1_R[30], U__d1, U__d0, P[68]);
  U4DPPG_31_19 U31 (P[70], O_R[69], IN1_R[31], U__d1, U__d0, P[69]);
  U4DPPG_32_19 U32 (P[71], O_R[70], IN1_R[32], U__d1, U__d0, P[70]);
  U4DPPG_33_19 U33 (P[72], O_R[71], IN1_R[33], U__d1, U__d0, P[71]);
  U4DPPG_34_19 U34 (P[73], O_R[72], IN1_R[34], U__d1, U__d0, P[72]);
  U4DPPG_35_19 U35 (P[74], O_R[73], IN1_R[35], U__d1, U__d0, P[73]);
  U4DPPG_36_19 U36 (P[75], O_R[74], IN1_R[36], U__d1, U__d0, P[74]);
  U4DPPG_37_19 U37 (P[76], O_R[75], IN1_R[37], U__d1, U__d0, P[75]);
  U4DPPG_38_19 U38 (P[77], O_R[76], IN1_R[38], U__d1, U__d0, P[76]);
  U4DPPG_39_19 U39 (P[78], O_R[77], IN1_R[39], U__d1, U__d0, P[77]);
  U4DPPG_40_19 U40 (P[79], O_R[78], IN1_R[40], U__d1, U__d0, P[78]);
  U4DPPG_41_19 U41 (P[80], O_R[79], IN1_R[41], U__d1, U__d0, P[79]);
  U4DPPG_42_19 U42 (P[81], O_R[80], IN1_R[42], U__d1, U__d0, P[80]);
  U4DPPG_43_19 U43 (P[82], O_R[81], IN1_R[43], U__d1, U__d0, P[81]);
  U4DPPG_44_19 U44 (P[83], O_R[82], IN1_R[44], U__d1, U__d0, P[82]);
  U4DPPG_45_19 U45 (P[84], O_R[83], IN1_R[45], U__d1, U__d0, P[83]);
  U4DPPG_46_19 U46 (P[85], O_R[84], IN1_R[46], U__d1, U__d0, P[84]);
  U4DPPG_47_19 U47 (P[86], O_R[85], IN1_R[47], U__d1, U__d0, P[85]);
  U4DPPG_48_19 U48 (P[87], O_R[86], IN1_R[48], U__d1, U__d0, P[86]);
  U4DPPG_49_19 U49 (P[88], O_R[87], IN1_R[49], U__d1, U__d0, P[87]);
  U4DPPG_50_19 U50 (P[89], O_R[88], IN1_R[50], U__d1, U__d0, P[88]);
  U4DPPG_51_19 U51 (P[90], O_R[89], IN1_R[51], U__d1, U__d0, P[89]);
  U4DPPG_52_19 U52 (P[91], O_R[90], IN1_R[52], U__d1, U__d0, P[90]);
  U4DPPG_53_19 U53 (P[92], O_R[91], IN1_R[53], U__d1, U__d0, P[91]);
  U4DPPG_54_19 U54 (P[93], O_R[92], IN1_R[54], U__d1, U__d0, P[92]);
  U4DPPG_55_19 U55 (P[94], O_R[93], IN1_R[55], U__d1, U__d0, P[93]);
  U4DPPG_56_19 U56 (P[95], O_R[94], IN1_R[56], U__d1, U__d0, P[94]);
  U4DPPG_57_19 U57 (P[96], O_R[95], IN1_R[57], U__d1, U__d0, P[95]);
  U4DPPG_58_19 U58 (P[97], O_R[96], IN1_R[58], U__d1, U__d0, P[96]);
  U4DPPG_59_19 U59 (P[98], O_R[97], IN1_R[59], U__d1, U__d0, P[97]);
  U4DPPG_60_19 U60 (P[99], O_R[98], IN1_R[60], U__d1, U__d0, P[98]);
  U4DPPG_61_19 U61 (P[100], O_R[99], IN1_R[61], U__d1, U__d0, P[99]);
  U4DPPG_62_19 U62 (P[101], O_R[100], IN1_R[62], U__d1, U__d0, P[100]);
  U4DPPGH_63_19 U63 (O_T, O_R[101], IN1_T, U__d1, U__d0, P[101]);
endmodule

module TCU4VPPG_63_0_2 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [67:4] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [67:5] P;
  U4DPPGL_0_2 U0 (P[5], O_R[4], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_2 U1 (P[6], O_R[5], IN1_R[1], U__d1, U__d0, P[5]);
  U4DPPG_2_2 U2 (P[7], O_R[6], IN1_R[2], U__d1, U__d0, P[6]);
  U4DPPG_3_2 U3 (P[8], O_R[7], IN1_R[3], U__d1, U__d0, P[7]);
  U4DPPG_4_2 U4 (P[9], O_R[8], IN1_R[4], U__d1, U__d0, P[8]);
  U4DPPG_5_2 U5 (P[10], O_R[9], IN1_R[5], U__d1, U__d0, P[9]);
  U4DPPG_6_2 U6 (P[11], O_R[10], IN1_R[6], U__d1, U__d0, P[10]);
  U4DPPG_7_2 U7 (P[12], O_R[11], IN1_R[7], U__d1, U__d0, P[11]);
  U4DPPG_8_2 U8 (P[13], O_R[12], IN1_R[8], U__d1, U__d0, P[12]);
  U4DPPG_9_2 U9 (P[14], O_R[13], IN1_R[9], U__d1, U__d0, P[13]);
  U4DPPG_10_2 U10 (P[15], O_R[14], IN1_R[10], U__d1, U__d0, P[14]);
  U4DPPG_11_2 U11 (P[16], O_R[15], IN1_R[11], U__d1, U__d0, P[15]);
  U4DPPG_12_2 U12 (P[17], O_R[16], IN1_R[12], U__d1, U__d0, P[16]);
  U4DPPG_13_2 U13 (P[18], O_R[17], IN1_R[13], U__d1, U__d0, P[17]);
  U4DPPG_14_2 U14 (P[19], O_R[18], IN1_R[14], U__d1, U__d0, P[18]);
  U4DPPG_15_2 U15 (P[20], O_R[19], IN1_R[15], U__d1, U__d0, P[19]);
  U4DPPG_16_2 U16 (P[21], O_R[20], IN1_R[16], U__d1, U__d0, P[20]);
  U4DPPG_17_2 U17 (P[22], O_R[21], IN1_R[17], U__d1, U__d0, P[21]);
  U4DPPG_18_2 U18 (P[23], O_R[22], IN1_R[18], U__d1, U__d0, P[22]);
  U4DPPG_19_2 U19 (P[24], O_R[23], IN1_R[19], U__d1, U__d0, P[23]);
  U4DPPG_20_2 U20 (P[25], O_R[24], IN1_R[20], U__d1, U__d0, P[24]);
  U4DPPG_21_2 U21 (P[26], O_R[25], IN1_R[21], U__d1, U__d0, P[25]);
  U4DPPG_22_2 U22 (P[27], O_R[26], IN1_R[22], U__d1, U__d0, P[26]);
  U4DPPG_23_2 U23 (P[28], O_R[27], IN1_R[23], U__d1, U__d0, P[27]);
  U4DPPG_24_2 U24 (P[29], O_R[28], IN1_R[24], U__d1, U__d0, P[28]);
  U4DPPG_25_2 U25 (P[30], O_R[29], IN1_R[25], U__d1, U__d0, P[29]);
  U4DPPG_26_2 U26 (P[31], O_R[30], IN1_R[26], U__d1, U__d0, P[30]);
  U4DPPG_27_2 U27 (P[32], O_R[31], IN1_R[27], U__d1, U__d0, P[31]);
  U4DPPG_28_2 U28 (P[33], O_R[32], IN1_R[28], U__d1, U__d0, P[32]);
  U4DPPG_29_2 U29 (P[34], O_R[33], IN1_R[29], U__d1, U__d0, P[33]);
  U4DPPG_30_2 U30 (P[35], O_R[34], IN1_R[30], U__d1, U__d0, P[34]);
  U4DPPG_31_2 U31 (P[36], O_R[35], IN1_R[31], U__d1, U__d0, P[35]);
  U4DPPG_32_2 U32 (P[37], O_R[36], IN1_R[32], U__d1, U__d0, P[36]);
  U4DPPG_33_2 U33 (P[38], O_R[37], IN1_R[33], U__d1, U__d0, P[37]);
  U4DPPG_34_2 U34 (P[39], O_R[38], IN1_R[34], U__d1, U__d0, P[38]);
  U4DPPG_35_2 U35 (P[40], O_R[39], IN1_R[35], U__d1, U__d0, P[39]);
  U4DPPG_36_2 U36 (P[41], O_R[40], IN1_R[36], U__d1, U__d0, P[40]);
  U4DPPG_37_2 U37 (P[42], O_R[41], IN1_R[37], U__d1, U__d0, P[41]);
  U4DPPG_38_2 U38 (P[43], O_R[42], IN1_R[38], U__d1, U__d0, P[42]);
  U4DPPG_39_2 U39 (P[44], O_R[43], IN1_R[39], U__d1, U__d0, P[43]);
  U4DPPG_40_2 U40 (P[45], O_R[44], IN1_R[40], U__d1, U__d0, P[44]);
  U4DPPG_41_2 U41 (P[46], O_R[45], IN1_R[41], U__d1, U__d0, P[45]);
  U4DPPG_42_2 U42 (P[47], O_R[46], IN1_R[42], U__d1, U__d0, P[46]);
  U4DPPG_43_2 U43 (P[48], O_R[47], IN1_R[43], U__d1, U__d0, P[47]);
  U4DPPG_44_2 U44 (P[49], O_R[48], IN1_R[44], U__d1, U__d0, P[48]);
  U4DPPG_45_2 U45 (P[50], O_R[49], IN1_R[45], U__d1, U__d0, P[49]);
  U4DPPG_46_2 U46 (P[51], O_R[50], IN1_R[46], U__d1, U__d0, P[50]);
  U4DPPG_47_2 U47 (P[52], O_R[51], IN1_R[47], U__d1, U__d0, P[51]);
  U4DPPG_48_2 U48 (P[53], O_R[52], IN1_R[48], U__d1, U__d0, P[52]);
  U4DPPG_49_2 U49 (P[54], O_R[53], IN1_R[49], U__d1, U__d0, P[53]);
  U4DPPG_50_2 U50 (P[55], O_R[54], IN1_R[50], U__d1, U__d0, P[54]);
  U4DPPG_51_2 U51 (P[56], O_R[55], IN1_R[51], U__d1, U__d0, P[55]);
  U4DPPG_52_2 U52 (P[57], O_R[56], IN1_R[52], U__d1, U__d0, P[56]);
  U4DPPG_53_2 U53 (P[58], O_R[57], IN1_R[53], U__d1, U__d0, P[57]);
  U4DPPG_54_2 U54 (P[59], O_R[58], IN1_R[54], U__d1, U__d0, P[58]);
  U4DPPG_55_2 U55 (P[60], O_R[59], IN1_R[55], U__d1, U__d0, P[59]);
  U4DPPG_56_2 U56 (P[61], O_R[60], IN1_R[56], U__d1, U__d0, P[60]);
  U4DPPG_57_2 U57 (P[62], O_R[61], IN1_R[57], U__d1, U__d0, P[61]);
  U4DPPG_58_2 U58 (P[63], O_R[62], IN1_R[58], U__d1, U__d0, P[62]);
  U4DPPG_59_2 U59 (P[64], O_R[63], IN1_R[59], U__d1, U__d0, P[63]);
  U4DPPG_60_2 U60 (P[65], O_R[64], IN1_R[60], U__d1, U__d0, P[64]);
  U4DPPG_61_2 U61 (P[66], O_R[65], IN1_R[61], U__d1, U__d0, P[65]);
  U4DPPG_62_2 U62 (P[67], O_R[66], IN1_R[62], U__d1, U__d0, P[66]);
  U4DPPGH_63_2 U63 (O_T, O_R[67], IN1_T, U__d1, U__d0, P[67]);
endmodule

module TCU4VPPG_63_0_20 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [103:40] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [103:41] P;
  U4DPPGL_0_20 U0 (P[41], O_R[40], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_20 U1 (P[42], O_R[41], IN1_R[1], U__d1, U__d0, P[41]);
  U4DPPG_2_20 U2 (P[43], O_R[42], IN1_R[2], U__d1, U__d0, P[42]);
  U4DPPG_3_20 U3 (P[44], O_R[43], IN1_R[3], U__d1, U__d0, P[43]);
  U4DPPG_4_20 U4 (P[45], O_R[44], IN1_R[4], U__d1, U__d0, P[44]);
  U4DPPG_5_20 U5 (P[46], O_R[45], IN1_R[5], U__d1, U__d0, P[45]);
  U4DPPG_6_20 U6 (P[47], O_R[46], IN1_R[6], U__d1, U__d0, P[46]);
  U4DPPG_7_20 U7 (P[48], O_R[47], IN1_R[7], U__d1, U__d0, P[47]);
  U4DPPG_8_20 U8 (P[49], O_R[48], IN1_R[8], U__d1, U__d0, P[48]);
  U4DPPG_9_20 U9 (P[50], O_R[49], IN1_R[9], U__d1, U__d0, P[49]);
  U4DPPG_10_20 U10 (P[51], O_R[50], IN1_R[10], U__d1, U__d0, P[50]);
  U4DPPG_11_20 U11 (P[52], O_R[51], IN1_R[11], U__d1, U__d0, P[51]);
  U4DPPG_12_20 U12 (P[53], O_R[52], IN1_R[12], U__d1, U__d0, P[52]);
  U4DPPG_13_20 U13 (P[54], O_R[53], IN1_R[13], U__d1, U__d0, P[53]);
  U4DPPG_14_20 U14 (P[55], O_R[54], IN1_R[14], U__d1, U__d0, P[54]);
  U4DPPG_15_20 U15 (P[56], O_R[55], IN1_R[15], U__d1, U__d0, P[55]);
  U4DPPG_16_20 U16 (P[57], O_R[56], IN1_R[16], U__d1, U__d0, P[56]);
  U4DPPG_17_20 U17 (P[58], O_R[57], IN1_R[17], U__d1, U__d0, P[57]);
  U4DPPG_18_20 U18 (P[59], O_R[58], IN1_R[18], U__d1, U__d0, P[58]);
  U4DPPG_19_20 U19 (P[60], O_R[59], IN1_R[19], U__d1, U__d0, P[59]);
  U4DPPG_20_20 U20 (P[61], O_R[60], IN1_R[20], U__d1, U__d0, P[60]);
  U4DPPG_21_20 U21 (P[62], O_R[61], IN1_R[21], U__d1, U__d0, P[61]);
  U4DPPG_22_20 U22 (P[63], O_R[62], IN1_R[22], U__d1, U__d0, P[62]);
  U4DPPG_23_20 U23 (P[64], O_R[63], IN1_R[23], U__d1, U__d0, P[63]);
  U4DPPG_24_20 U24 (P[65], O_R[64], IN1_R[24], U__d1, U__d0, P[64]);
  U4DPPG_25_20 U25 (P[66], O_R[65], IN1_R[25], U__d1, U__d0, P[65]);
  U4DPPG_26_20 U26 (P[67], O_R[66], IN1_R[26], U__d1, U__d0, P[66]);
  U4DPPG_27_20 U27 (P[68], O_R[67], IN1_R[27], U__d1, U__d0, P[67]);
  U4DPPG_28_20 U28 (P[69], O_R[68], IN1_R[28], U__d1, U__d0, P[68]);
  U4DPPG_29_20 U29 (P[70], O_R[69], IN1_R[29], U__d1, U__d0, P[69]);
  U4DPPG_30_20 U30 (P[71], O_R[70], IN1_R[30], U__d1, U__d0, P[70]);
  U4DPPG_31_20 U31 (P[72], O_R[71], IN1_R[31], U__d1, U__d0, P[71]);
  U4DPPG_32_20 U32 (P[73], O_R[72], IN1_R[32], U__d1, U__d0, P[72]);
  U4DPPG_33_20 U33 (P[74], O_R[73], IN1_R[33], U__d1, U__d0, P[73]);
  U4DPPG_34_20 U34 (P[75], O_R[74], IN1_R[34], U__d1, U__d0, P[74]);
  U4DPPG_35_20 U35 (P[76], O_R[75], IN1_R[35], U__d1, U__d0, P[75]);
  U4DPPG_36_20 U36 (P[77], O_R[76], IN1_R[36], U__d1, U__d0, P[76]);
  U4DPPG_37_20 U37 (P[78], O_R[77], IN1_R[37], U__d1, U__d0, P[77]);
  U4DPPG_38_20 U38 (P[79], O_R[78], IN1_R[38], U__d1, U__d0, P[78]);
  U4DPPG_39_20 U39 (P[80], O_R[79], IN1_R[39], U__d1, U__d0, P[79]);
  U4DPPG_40_20 U40 (P[81], O_R[80], IN1_R[40], U__d1, U__d0, P[80]);
  U4DPPG_41_20 U41 (P[82], O_R[81], IN1_R[41], U__d1, U__d0, P[81]);
  U4DPPG_42_20 U42 (P[83], O_R[82], IN1_R[42], U__d1, U__d0, P[82]);
  U4DPPG_43_20 U43 (P[84], O_R[83], IN1_R[43], U__d1, U__d0, P[83]);
  U4DPPG_44_20 U44 (P[85], O_R[84], IN1_R[44], U__d1, U__d0, P[84]);
  U4DPPG_45_20 U45 (P[86], O_R[85], IN1_R[45], U__d1, U__d0, P[85]);
  U4DPPG_46_20 U46 (P[87], O_R[86], IN1_R[46], U__d1, U__d0, P[86]);
  U4DPPG_47_20 U47 (P[88], O_R[87], IN1_R[47], U__d1, U__d0, P[87]);
  U4DPPG_48_20 U48 (P[89], O_R[88], IN1_R[48], U__d1, U__d0, P[88]);
  U4DPPG_49_20 U49 (P[90], O_R[89], IN1_R[49], U__d1, U__d0, P[89]);
  U4DPPG_50_20 U50 (P[91], O_R[90], IN1_R[50], U__d1, U__d0, P[90]);
  U4DPPG_51_20 U51 (P[92], O_R[91], IN1_R[51], U__d1, U__d0, P[91]);
  U4DPPG_52_20 U52 (P[93], O_R[92], IN1_R[52], U__d1, U__d0, P[92]);
  U4DPPG_53_20 U53 (P[94], O_R[93], IN1_R[53], U__d1, U__d0, P[93]);
  U4DPPG_54_20 U54 (P[95], O_R[94], IN1_R[54], U__d1, U__d0, P[94]);
  U4DPPG_55_20 U55 (P[96], O_R[95], IN1_R[55], U__d1, U__d0, P[95]);
  U4DPPG_56_20 U56 (P[97], O_R[96], IN1_R[56], U__d1, U__d0, P[96]);
  U4DPPG_57_20 U57 (P[98], O_R[97], IN1_R[57], U__d1, U__d0, P[97]);
  U4DPPG_58_20 U58 (P[99], O_R[98], IN1_R[58], U__d1, U__d0, P[98]);
  U4DPPG_59_20 U59 (P[100], O_R[99], IN1_R[59], U__d1, U__d0, P[99]);
  U4DPPG_60_20 U60 (P[101], O_R[100], IN1_R[60], U__d1, U__d0, P[100]);
  U4DPPG_61_20 U61 (P[102], O_R[101], IN1_R[61], U__d1, U__d0, P[101]);
  U4DPPG_62_20 U62 (P[103], O_R[102], IN1_R[62], U__d1, U__d0, P[102]);
  U4DPPGH_63_20 U63 (O_T, O_R[103], IN1_T, U__d1, U__d0, P[103]);
endmodule

module TCU4VPPG_63_0_21 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [105:42] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [105:43] P;
  U4DPPGL_0_21 U0 (P[43], O_R[42], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_21 U1 (P[44], O_R[43], IN1_R[1], U__d1, U__d0, P[43]);
  U4DPPG_2_21 U2 (P[45], O_R[44], IN1_R[2], U__d1, U__d0, P[44]);
  U4DPPG_3_21 U3 (P[46], O_R[45], IN1_R[3], U__d1, U__d0, P[45]);
  U4DPPG_4_21 U4 (P[47], O_R[46], IN1_R[4], U__d1, U__d0, P[46]);
  U4DPPG_5_21 U5 (P[48], O_R[47], IN1_R[5], U__d1, U__d0, P[47]);
  U4DPPG_6_21 U6 (P[49], O_R[48], IN1_R[6], U__d1, U__d0, P[48]);
  U4DPPG_7_21 U7 (P[50], O_R[49], IN1_R[7], U__d1, U__d0, P[49]);
  U4DPPG_8_21 U8 (P[51], O_R[50], IN1_R[8], U__d1, U__d0, P[50]);
  U4DPPG_9_21 U9 (P[52], O_R[51], IN1_R[9], U__d1, U__d0, P[51]);
  U4DPPG_10_21 U10 (P[53], O_R[52], IN1_R[10], U__d1, U__d0, P[52]);
  U4DPPG_11_21 U11 (P[54], O_R[53], IN1_R[11], U__d1, U__d0, P[53]);
  U4DPPG_12_21 U12 (P[55], O_R[54], IN1_R[12], U__d1, U__d0, P[54]);
  U4DPPG_13_21 U13 (P[56], O_R[55], IN1_R[13], U__d1, U__d0, P[55]);
  U4DPPG_14_21 U14 (P[57], O_R[56], IN1_R[14], U__d1, U__d0, P[56]);
  U4DPPG_15_21 U15 (P[58], O_R[57], IN1_R[15], U__d1, U__d0, P[57]);
  U4DPPG_16_21 U16 (P[59], O_R[58], IN1_R[16], U__d1, U__d0, P[58]);
  U4DPPG_17_21 U17 (P[60], O_R[59], IN1_R[17], U__d1, U__d0, P[59]);
  U4DPPG_18_21 U18 (P[61], O_R[60], IN1_R[18], U__d1, U__d0, P[60]);
  U4DPPG_19_21 U19 (P[62], O_R[61], IN1_R[19], U__d1, U__d0, P[61]);
  U4DPPG_20_21 U20 (P[63], O_R[62], IN1_R[20], U__d1, U__d0, P[62]);
  U4DPPG_21_21 U21 (P[64], O_R[63], IN1_R[21], U__d1, U__d0, P[63]);
  U4DPPG_22_21 U22 (P[65], O_R[64], IN1_R[22], U__d1, U__d0, P[64]);
  U4DPPG_23_21 U23 (P[66], O_R[65], IN1_R[23], U__d1, U__d0, P[65]);
  U4DPPG_24_21 U24 (P[67], O_R[66], IN1_R[24], U__d1, U__d0, P[66]);
  U4DPPG_25_21 U25 (P[68], O_R[67], IN1_R[25], U__d1, U__d0, P[67]);
  U4DPPG_26_21 U26 (P[69], O_R[68], IN1_R[26], U__d1, U__d0, P[68]);
  U4DPPG_27_21 U27 (P[70], O_R[69], IN1_R[27], U__d1, U__d0, P[69]);
  U4DPPG_28_21 U28 (P[71], O_R[70], IN1_R[28], U__d1, U__d0, P[70]);
  U4DPPG_29_21 U29 (P[72], O_R[71], IN1_R[29], U__d1, U__d0, P[71]);
  U4DPPG_30_21 U30 (P[73], O_R[72], IN1_R[30], U__d1, U__d0, P[72]);
  U4DPPG_31_21 U31 (P[74], O_R[73], IN1_R[31], U__d1, U__d0, P[73]);
  U4DPPG_32_21 U32 (P[75], O_R[74], IN1_R[32], U__d1, U__d0, P[74]);
  U4DPPG_33_21 U33 (P[76], O_R[75], IN1_R[33], U__d1, U__d0, P[75]);
  U4DPPG_34_21 U34 (P[77], O_R[76], IN1_R[34], U__d1, U__d0, P[76]);
  U4DPPG_35_21 U35 (P[78], O_R[77], IN1_R[35], U__d1, U__d0, P[77]);
  U4DPPG_36_21 U36 (P[79], O_R[78], IN1_R[36], U__d1, U__d0, P[78]);
  U4DPPG_37_21 U37 (P[80], O_R[79], IN1_R[37], U__d1, U__d0, P[79]);
  U4DPPG_38_21 U38 (P[81], O_R[80], IN1_R[38], U__d1, U__d0, P[80]);
  U4DPPG_39_21 U39 (P[82], O_R[81], IN1_R[39], U__d1, U__d0, P[81]);
  U4DPPG_40_21 U40 (P[83], O_R[82], IN1_R[40], U__d1, U__d0, P[82]);
  U4DPPG_41_21 U41 (P[84], O_R[83], IN1_R[41], U__d1, U__d0, P[83]);
  U4DPPG_42_21 U42 (P[85], O_R[84], IN1_R[42], U__d1, U__d0, P[84]);
  U4DPPG_43_21 U43 (P[86], O_R[85], IN1_R[43], U__d1, U__d0, P[85]);
  U4DPPG_44_21 U44 (P[87], O_R[86], IN1_R[44], U__d1, U__d0, P[86]);
  U4DPPG_45_21 U45 (P[88], O_R[87], IN1_R[45], U__d1, U__d0, P[87]);
  U4DPPG_46_21 U46 (P[89], O_R[88], IN1_R[46], U__d1, U__d0, P[88]);
  U4DPPG_47_21 U47 (P[90], O_R[89], IN1_R[47], U__d1, U__d0, P[89]);
  U4DPPG_48_21 U48 (P[91], O_R[90], IN1_R[48], U__d1, U__d0, P[90]);
  U4DPPG_49_21 U49 (P[92], O_R[91], IN1_R[49], U__d1, U__d0, P[91]);
  U4DPPG_50_21 U50 (P[93], O_R[92], IN1_R[50], U__d1, U__d0, P[92]);
  U4DPPG_51_21 U51 (P[94], O_R[93], IN1_R[51], U__d1, U__d0, P[93]);
  U4DPPG_52_21 U52 (P[95], O_R[94], IN1_R[52], U__d1, U__d0, P[94]);
  U4DPPG_53_21 U53 (P[96], O_R[95], IN1_R[53], U__d1, U__d0, P[95]);
  U4DPPG_54_21 U54 (P[97], O_R[96], IN1_R[54], U__d1, U__d0, P[96]);
  U4DPPG_55_21 U55 (P[98], O_R[97], IN1_R[55], U__d1, U__d0, P[97]);
  U4DPPG_56_21 U56 (P[99], O_R[98], IN1_R[56], U__d1, U__d0, P[98]);
  U4DPPG_57_21 U57 (P[100], O_R[99], IN1_R[57], U__d1, U__d0, P[99]);
  U4DPPG_58_21 U58 (P[101], O_R[100], IN1_R[58], U__d1, U__d0, P[100]);
  U4DPPG_59_21 U59 (P[102], O_R[101], IN1_R[59], U__d1, U__d0, P[101]);
  U4DPPG_60_21 U60 (P[103], O_R[102], IN1_R[60], U__d1, U__d0, P[102]);
  U4DPPG_61_21 U61 (P[104], O_R[103], IN1_R[61], U__d1, U__d0, P[103]);
  U4DPPG_62_21 U62 (P[105], O_R[104], IN1_R[62], U__d1, U__d0, P[104]);
  U4DPPGH_63_21 U63 (O_T, O_R[105], IN1_T, U__d1, U__d0, P[105]);
endmodule

module TCU4VPPG_63_0_22 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [107:44] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [107:45] P;
  U4DPPGL_0_22 U0 (P[45], O_R[44], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_22 U1 (P[46], O_R[45], IN1_R[1], U__d1, U__d0, P[45]);
  U4DPPG_2_22 U2 (P[47], O_R[46], IN1_R[2], U__d1, U__d0, P[46]);
  U4DPPG_3_22 U3 (P[48], O_R[47], IN1_R[3], U__d1, U__d0, P[47]);
  U4DPPG_4_22 U4 (P[49], O_R[48], IN1_R[4], U__d1, U__d0, P[48]);
  U4DPPG_5_22 U5 (P[50], O_R[49], IN1_R[5], U__d1, U__d0, P[49]);
  U4DPPG_6_22 U6 (P[51], O_R[50], IN1_R[6], U__d1, U__d0, P[50]);
  U4DPPG_7_22 U7 (P[52], O_R[51], IN1_R[7], U__d1, U__d0, P[51]);
  U4DPPG_8_22 U8 (P[53], O_R[52], IN1_R[8], U__d1, U__d0, P[52]);
  U4DPPG_9_22 U9 (P[54], O_R[53], IN1_R[9], U__d1, U__d0, P[53]);
  U4DPPG_10_22 U10 (P[55], O_R[54], IN1_R[10], U__d1, U__d0, P[54]);
  U4DPPG_11_22 U11 (P[56], O_R[55], IN1_R[11], U__d1, U__d0, P[55]);
  U4DPPG_12_22 U12 (P[57], O_R[56], IN1_R[12], U__d1, U__d0, P[56]);
  U4DPPG_13_22 U13 (P[58], O_R[57], IN1_R[13], U__d1, U__d0, P[57]);
  U4DPPG_14_22 U14 (P[59], O_R[58], IN1_R[14], U__d1, U__d0, P[58]);
  U4DPPG_15_22 U15 (P[60], O_R[59], IN1_R[15], U__d1, U__d0, P[59]);
  U4DPPG_16_22 U16 (P[61], O_R[60], IN1_R[16], U__d1, U__d0, P[60]);
  U4DPPG_17_22 U17 (P[62], O_R[61], IN1_R[17], U__d1, U__d0, P[61]);
  U4DPPG_18_22 U18 (P[63], O_R[62], IN1_R[18], U__d1, U__d0, P[62]);
  U4DPPG_19_22 U19 (P[64], O_R[63], IN1_R[19], U__d1, U__d0, P[63]);
  U4DPPG_20_22 U20 (P[65], O_R[64], IN1_R[20], U__d1, U__d0, P[64]);
  U4DPPG_21_22 U21 (P[66], O_R[65], IN1_R[21], U__d1, U__d0, P[65]);
  U4DPPG_22_22 U22 (P[67], O_R[66], IN1_R[22], U__d1, U__d0, P[66]);
  U4DPPG_23_22 U23 (P[68], O_R[67], IN1_R[23], U__d1, U__d0, P[67]);
  U4DPPG_24_22 U24 (P[69], O_R[68], IN1_R[24], U__d1, U__d0, P[68]);
  U4DPPG_25_22 U25 (P[70], O_R[69], IN1_R[25], U__d1, U__d0, P[69]);
  U4DPPG_26_22 U26 (P[71], O_R[70], IN1_R[26], U__d1, U__d0, P[70]);
  U4DPPG_27_22 U27 (P[72], O_R[71], IN1_R[27], U__d1, U__d0, P[71]);
  U4DPPG_28_22 U28 (P[73], O_R[72], IN1_R[28], U__d1, U__d0, P[72]);
  U4DPPG_29_22 U29 (P[74], O_R[73], IN1_R[29], U__d1, U__d0, P[73]);
  U4DPPG_30_22 U30 (P[75], O_R[74], IN1_R[30], U__d1, U__d0, P[74]);
  U4DPPG_31_22 U31 (P[76], O_R[75], IN1_R[31], U__d1, U__d0, P[75]);
  U4DPPG_32_22 U32 (P[77], O_R[76], IN1_R[32], U__d1, U__d0, P[76]);
  U4DPPG_33_22 U33 (P[78], O_R[77], IN1_R[33], U__d1, U__d0, P[77]);
  U4DPPG_34_22 U34 (P[79], O_R[78], IN1_R[34], U__d1, U__d0, P[78]);
  U4DPPG_35_22 U35 (P[80], O_R[79], IN1_R[35], U__d1, U__d0, P[79]);
  U4DPPG_36_22 U36 (P[81], O_R[80], IN1_R[36], U__d1, U__d0, P[80]);
  U4DPPG_37_22 U37 (P[82], O_R[81], IN1_R[37], U__d1, U__d0, P[81]);
  U4DPPG_38_22 U38 (P[83], O_R[82], IN1_R[38], U__d1, U__d0, P[82]);
  U4DPPG_39_22 U39 (P[84], O_R[83], IN1_R[39], U__d1, U__d0, P[83]);
  U4DPPG_40_22 U40 (P[85], O_R[84], IN1_R[40], U__d1, U__d0, P[84]);
  U4DPPG_41_22 U41 (P[86], O_R[85], IN1_R[41], U__d1, U__d0, P[85]);
  U4DPPG_42_22 U42 (P[87], O_R[86], IN1_R[42], U__d1, U__d0, P[86]);
  U4DPPG_43_22 U43 (P[88], O_R[87], IN1_R[43], U__d1, U__d0, P[87]);
  U4DPPG_44_22 U44 (P[89], O_R[88], IN1_R[44], U__d1, U__d0, P[88]);
  U4DPPG_45_22 U45 (P[90], O_R[89], IN1_R[45], U__d1, U__d0, P[89]);
  U4DPPG_46_22 U46 (P[91], O_R[90], IN1_R[46], U__d1, U__d0, P[90]);
  U4DPPG_47_22 U47 (P[92], O_R[91], IN1_R[47], U__d1, U__d0, P[91]);
  U4DPPG_48_22 U48 (P[93], O_R[92], IN1_R[48], U__d1, U__d0, P[92]);
  U4DPPG_49_22 U49 (P[94], O_R[93], IN1_R[49], U__d1, U__d0, P[93]);
  U4DPPG_50_22 U50 (P[95], O_R[94], IN1_R[50], U__d1, U__d0, P[94]);
  U4DPPG_51_22 U51 (P[96], O_R[95], IN1_R[51], U__d1, U__d0, P[95]);
  U4DPPG_52_22 U52 (P[97], O_R[96], IN1_R[52], U__d1, U__d0, P[96]);
  U4DPPG_53_22 U53 (P[98], O_R[97], IN1_R[53], U__d1, U__d0, P[97]);
  U4DPPG_54_22 U54 (P[99], O_R[98], IN1_R[54], U__d1, U__d0, P[98]);
  U4DPPG_55_22 U55 (P[100], O_R[99], IN1_R[55], U__d1, U__d0, P[99]);
  U4DPPG_56_22 U56 (P[101], O_R[100], IN1_R[56], U__d1, U__d0, P[100]);
  U4DPPG_57_22 U57 (P[102], O_R[101], IN1_R[57], U__d1, U__d0, P[101]);
  U4DPPG_58_22 U58 (P[103], O_R[102], IN1_R[58], U__d1, U__d0, P[102]);
  U4DPPG_59_22 U59 (P[104], O_R[103], IN1_R[59], U__d1, U__d0, P[103]);
  U4DPPG_60_22 U60 (P[105], O_R[104], IN1_R[60], U__d1, U__d0, P[104]);
  U4DPPG_61_22 U61 (P[106], O_R[105], IN1_R[61], U__d1, U__d0, P[105]);
  U4DPPG_62_22 U62 (P[107], O_R[106], IN1_R[62], U__d1, U__d0, P[106]);
  U4DPPGH_63_22 U63 (O_T, O_R[107], IN1_T, U__d1, U__d0, P[107]);
endmodule

module TCU4VPPG_63_0_23 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [109:46] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [109:47] P;
  U4DPPGL_0_23 U0 (P[47], O_R[46], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_23 U1 (P[48], O_R[47], IN1_R[1], U__d1, U__d0, P[47]);
  U4DPPG_2_23 U2 (P[49], O_R[48], IN1_R[2], U__d1, U__d0, P[48]);
  U4DPPG_3_23 U3 (P[50], O_R[49], IN1_R[3], U__d1, U__d0, P[49]);
  U4DPPG_4_23 U4 (P[51], O_R[50], IN1_R[4], U__d1, U__d0, P[50]);
  U4DPPG_5_23 U5 (P[52], O_R[51], IN1_R[5], U__d1, U__d0, P[51]);
  U4DPPG_6_23 U6 (P[53], O_R[52], IN1_R[6], U__d1, U__d0, P[52]);
  U4DPPG_7_23 U7 (P[54], O_R[53], IN1_R[7], U__d1, U__d0, P[53]);
  U4DPPG_8_23 U8 (P[55], O_R[54], IN1_R[8], U__d1, U__d0, P[54]);
  U4DPPG_9_23 U9 (P[56], O_R[55], IN1_R[9], U__d1, U__d0, P[55]);
  U4DPPG_10_23 U10 (P[57], O_R[56], IN1_R[10], U__d1, U__d0, P[56]);
  U4DPPG_11_23 U11 (P[58], O_R[57], IN1_R[11], U__d1, U__d0, P[57]);
  U4DPPG_12_23 U12 (P[59], O_R[58], IN1_R[12], U__d1, U__d0, P[58]);
  U4DPPG_13_23 U13 (P[60], O_R[59], IN1_R[13], U__d1, U__d0, P[59]);
  U4DPPG_14_23 U14 (P[61], O_R[60], IN1_R[14], U__d1, U__d0, P[60]);
  U4DPPG_15_23 U15 (P[62], O_R[61], IN1_R[15], U__d1, U__d0, P[61]);
  U4DPPG_16_23 U16 (P[63], O_R[62], IN1_R[16], U__d1, U__d0, P[62]);
  U4DPPG_17_23 U17 (P[64], O_R[63], IN1_R[17], U__d1, U__d0, P[63]);
  U4DPPG_18_23 U18 (P[65], O_R[64], IN1_R[18], U__d1, U__d0, P[64]);
  U4DPPG_19_23 U19 (P[66], O_R[65], IN1_R[19], U__d1, U__d0, P[65]);
  U4DPPG_20_23 U20 (P[67], O_R[66], IN1_R[20], U__d1, U__d0, P[66]);
  U4DPPG_21_23 U21 (P[68], O_R[67], IN1_R[21], U__d1, U__d0, P[67]);
  U4DPPG_22_23 U22 (P[69], O_R[68], IN1_R[22], U__d1, U__d0, P[68]);
  U4DPPG_23_23 U23 (P[70], O_R[69], IN1_R[23], U__d1, U__d0, P[69]);
  U4DPPG_24_23 U24 (P[71], O_R[70], IN1_R[24], U__d1, U__d0, P[70]);
  U4DPPG_25_23 U25 (P[72], O_R[71], IN1_R[25], U__d1, U__d0, P[71]);
  U4DPPG_26_23 U26 (P[73], O_R[72], IN1_R[26], U__d1, U__d0, P[72]);
  U4DPPG_27_23 U27 (P[74], O_R[73], IN1_R[27], U__d1, U__d0, P[73]);
  U4DPPG_28_23 U28 (P[75], O_R[74], IN1_R[28], U__d1, U__d0, P[74]);
  U4DPPG_29_23 U29 (P[76], O_R[75], IN1_R[29], U__d1, U__d0, P[75]);
  U4DPPG_30_23 U30 (P[77], O_R[76], IN1_R[30], U__d1, U__d0, P[76]);
  U4DPPG_31_23 U31 (P[78], O_R[77], IN1_R[31], U__d1, U__d0, P[77]);
  U4DPPG_32_23 U32 (P[79], O_R[78], IN1_R[32], U__d1, U__d0, P[78]);
  U4DPPG_33_23 U33 (P[80], O_R[79], IN1_R[33], U__d1, U__d0, P[79]);
  U4DPPG_34_23 U34 (P[81], O_R[80], IN1_R[34], U__d1, U__d0, P[80]);
  U4DPPG_35_23 U35 (P[82], O_R[81], IN1_R[35], U__d1, U__d0, P[81]);
  U4DPPG_36_23 U36 (P[83], O_R[82], IN1_R[36], U__d1, U__d0, P[82]);
  U4DPPG_37_23 U37 (P[84], O_R[83], IN1_R[37], U__d1, U__d0, P[83]);
  U4DPPG_38_23 U38 (P[85], O_R[84], IN1_R[38], U__d1, U__d0, P[84]);
  U4DPPG_39_23 U39 (P[86], O_R[85], IN1_R[39], U__d1, U__d0, P[85]);
  U4DPPG_40_23 U40 (P[87], O_R[86], IN1_R[40], U__d1, U__d0, P[86]);
  U4DPPG_41_23 U41 (P[88], O_R[87], IN1_R[41], U__d1, U__d0, P[87]);
  U4DPPG_42_23 U42 (P[89], O_R[88], IN1_R[42], U__d1, U__d0, P[88]);
  U4DPPG_43_23 U43 (P[90], O_R[89], IN1_R[43], U__d1, U__d0, P[89]);
  U4DPPG_44_23 U44 (P[91], O_R[90], IN1_R[44], U__d1, U__d0, P[90]);
  U4DPPG_45_23 U45 (P[92], O_R[91], IN1_R[45], U__d1, U__d0, P[91]);
  U4DPPG_46_23 U46 (P[93], O_R[92], IN1_R[46], U__d1, U__d0, P[92]);
  U4DPPG_47_23 U47 (P[94], O_R[93], IN1_R[47], U__d1, U__d0, P[93]);
  U4DPPG_48_23 U48 (P[95], O_R[94], IN1_R[48], U__d1, U__d0, P[94]);
  U4DPPG_49_23 U49 (P[96], O_R[95], IN1_R[49], U__d1, U__d0, P[95]);
  U4DPPG_50_23 U50 (P[97], O_R[96], IN1_R[50], U__d1, U__d0, P[96]);
  U4DPPG_51_23 U51 (P[98], O_R[97], IN1_R[51], U__d1, U__d0, P[97]);
  U4DPPG_52_23 U52 (P[99], O_R[98], IN1_R[52], U__d1, U__d0, P[98]);
  U4DPPG_53_23 U53 (P[100], O_R[99], IN1_R[53], U__d1, U__d0, P[99]);
  U4DPPG_54_23 U54 (P[101], O_R[100], IN1_R[54], U__d1, U__d0, P[100]);
  U4DPPG_55_23 U55 (P[102], O_R[101], IN1_R[55], U__d1, U__d0, P[101]);
  U4DPPG_56_23 U56 (P[103], O_R[102], IN1_R[56], U__d1, U__d0, P[102]);
  U4DPPG_57_23 U57 (P[104], O_R[103], IN1_R[57], U__d1, U__d0, P[103]);
  U4DPPG_58_23 U58 (P[105], O_R[104], IN1_R[58], U__d1, U__d0, P[104]);
  U4DPPG_59_23 U59 (P[106], O_R[105], IN1_R[59], U__d1, U__d0, P[105]);
  U4DPPG_60_23 U60 (P[107], O_R[106], IN1_R[60], U__d1, U__d0, P[106]);
  U4DPPG_61_23 U61 (P[108], O_R[107], IN1_R[61], U__d1, U__d0, P[107]);
  U4DPPG_62_23 U62 (P[109], O_R[108], IN1_R[62], U__d1, U__d0, P[108]);
  U4DPPGH_63_23 U63 (O_T, O_R[109], IN1_T, U__d1, U__d0, P[109]);
endmodule

module TCU4VPPG_63_0_24 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [111:48] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [111:49] P;
  U4DPPGL_0_24 U0 (P[49], O_R[48], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_24 U1 (P[50], O_R[49], IN1_R[1], U__d1, U__d0, P[49]);
  U4DPPG_2_24 U2 (P[51], O_R[50], IN1_R[2], U__d1, U__d0, P[50]);
  U4DPPG_3_24 U3 (P[52], O_R[51], IN1_R[3], U__d1, U__d0, P[51]);
  U4DPPG_4_24 U4 (P[53], O_R[52], IN1_R[4], U__d1, U__d0, P[52]);
  U4DPPG_5_24 U5 (P[54], O_R[53], IN1_R[5], U__d1, U__d0, P[53]);
  U4DPPG_6_24 U6 (P[55], O_R[54], IN1_R[6], U__d1, U__d0, P[54]);
  U4DPPG_7_24 U7 (P[56], O_R[55], IN1_R[7], U__d1, U__d0, P[55]);
  U4DPPG_8_24 U8 (P[57], O_R[56], IN1_R[8], U__d1, U__d0, P[56]);
  U4DPPG_9_24 U9 (P[58], O_R[57], IN1_R[9], U__d1, U__d0, P[57]);
  U4DPPG_10_24 U10 (P[59], O_R[58], IN1_R[10], U__d1, U__d0, P[58]);
  U4DPPG_11_24 U11 (P[60], O_R[59], IN1_R[11], U__d1, U__d0, P[59]);
  U4DPPG_12_24 U12 (P[61], O_R[60], IN1_R[12], U__d1, U__d0, P[60]);
  U4DPPG_13_24 U13 (P[62], O_R[61], IN1_R[13], U__d1, U__d0, P[61]);
  U4DPPG_14_24 U14 (P[63], O_R[62], IN1_R[14], U__d1, U__d0, P[62]);
  U4DPPG_15_24 U15 (P[64], O_R[63], IN1_R[15], U__d1, U__d0, P[63]);
  U4DPPG_16_24 U16 (P[65], O_R[64], IN1_R[16], U__d1, U__d0, P[64]);
  U4DPPG_17_24 U17 (P[66], O_R[65], IN1_R[17], U__d1, U__d0, P[65]);
  U4DPPG_18_24 U18 (P[67], O_R[66], IN1_R[18], U__d1, U__d0, P[66]);
  U4DPPG_19_24 U19 (P[68], O_R[67], IN1_R[19], U__d1, U__d0, P[67]);
  U4DPPG_20_24 U20 (P[69], O_R[68], IN1_R[20], U__d1, U__d0, P[68]);
  U4DPPG_21_24 U21 (P[70], O_R[69], IN1_R[21], U__d1, U__d0, P[69]);
  U4DPPG_22_24 U22 (P[71], O_R[70], IN1_R[22], U__d1, U__d0, P[70]);
  U4DPPG_23_24 U23 (P[72], O_R[71], IN1_R[23], U__d1, U__d0, P[71]);
  U4DPPG_24_24 U24 (P[73], O_R[72], IN1_R[24], U__d1, U__d0, P[72]);
  U4DPPG_25_24 U25 (P[74], O_R[73], IN1_R[25], U__d1, U__d0, P[73]);
  U4DPPG_26_24 U26 (P[75], O_R[74], IN1_R[26], U__d1, U__d0, P[74]);
  U4DPPG_27_24 U27 (P[76], O_R[75], IN1_R[27], U__d1, U__d0, P[75]);
  U4DPPG_28_24 U28 (P[77], O_R[76], IN1_R[28], U__d1, U__d0, P[76]);
  U4DPPG_29_24 U29 (P[78], O_R[77], IN1_R[29], U__d1, U__d0, P[77]);
  U4DPPG_30_24 U30 (P[79], O_R[78], IN1_R[30], U__d1, U__d0, P[78]);
  U4DPPG_31_24 U31 (P[80], O_R[79], IN1_R[31], U__d1, U__d0, P[79]);
  U4DPPG_32_24 U32 (P[81], O_R[80], IN1_R[32], U__d1, U__d0, P[80]);
  U4DPPG_33_24 U33 (P[82], O_R[81], IN1_R[33], U__d1, U__d0, P[81]);
  U4DPPG_34_24 U34 (P[83], O_R[82], IN1_R[34], U__d1, U__d0, P[82]);
  U4DPPG_35_24 U35 (P[84], O_R[83], IN1_R[35], U__d1, U__d0, P[83]);
  U4DPPG_36_24 U36 (P[85], O_R[84], IN1_R[36], U__d1, U__d0, P[84]);
  U4DPPG_37_24 U37 (P[86], O_R[85], IN1_R[37], U__d1, U__d0, P[85]);
  U4DPPG_38_24 U38 (P[87], O_R[86], IN1_R[38], U__d1, U__d0, P[86]);
  U4DPPG_39_24 U39 (P[88], O_R[87], IN1_R[39], U__d1, U__d0, P[87]);
  U4DPPG_40_24 U40 (P[89], O_R[88], IN1_R[40], U__d1, U__d0, P[88]);
  U4DPPG_41_24 U41 (P[90], O_R[89], IN1_R[41], U__d1, U__d0, P[89]);
  U4DPPG_42_24 U42 (P[91], O_R[90], IN1_R[42], U__d1, U__d0, P[90]);
  U4DPPG_43_24 U43 (P[92], O_R[91], IN1_R[43], U__d1, U__d0, P[91]);
  U4DPPG_44_24 U44 (P[93], O_R[92], IN1_R[44], U__d1, U__d0, P[92]);
  U4DPPG_45_24 U45 (P[94], O_R[93], IN1_R[45], U__d1, U__d0, P[93]);
  U4DPPG_46_24 U46 (P[95], O_R[94], IN1_R[46], U__d1, U__d0, P[94]);
  U4DPPG_47_24 U47 (P[96], O_R[95], IN1_R[47], U__d1, U__d0, P[95]);
  U4DPPG_48_24 U48 (P[97], O_R[96], IN1_R[48], U__d1, U__d0, P[96]);
  U4DPPG_49_24 U49 (P[98], O_R[97], IN1_R[49], U__d1, U__d0, P[97]);
  U4DPPG_50_24 U50 (P[99], O_R[98], IN1_R[50], U__d1, U__d0, P[98]);
  U4DPPG_51_24 U51 (P[100], O_R[99], IN1_R[51], U__d1, U__d0, P[99]);
  U4DPPG_52_24 U52 (P[101], O_R[100], IN1_R[52], U__d1, U__d0, P[100]);
  U4DPPG_53_24 U53 (P[102], O_R[101], IN1_R[53], U__d1, U__d0, P[101]);
  U4DPPG_54_24 U54 (P[103], O_R[102], IN1_R[54], U__d1, U__d0, P[102]);
  U4DPPG_55_24 U55 (P[104], O_R[103], IN1_R[55], U__d1, U__d0, P[103]);
  U4DPPG_56_24 U56 (P[105], O_R[104], IN1_R[56], U__d1, U__d0, P[104]);
  U4DPPG_57_24 U57 (P[106], O_R[105], IN1_R[57], U__d1, U__d0, P[105]);
  U4DPPG_58_24 U58 (P[107], O_R[106], IN1_R[58], U__d1, U__d0, P[106]);
  U4DPPG_59_24 U59 (P[108], O_R[107], IN1_R[59], U__d1, U__d0, P[107]);
  U4DPPG_60_24 U60 (P[109], O_R[108], IN1_R[60], U__d1, U__d0, P[108]);
  U4DPPG_61_24 U61 (P[110], O_R[109], IN1_R[61], U__d1, U__d0, P[109]);
  U4DPPG_62_24 U62 (P[111], O_R[110], IN1_R[62], U__d1, U__d0, P[110]);
  U4DPPGH_63_24 U63 (O_T, O_R[111], IN1_T, U__d1, U__d0, P[111]);
endmodule

module TCU4VPPG_63_0_25 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [113:50] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [113:51] P;
  U4DPPGL_0_25 U0 (P[51], O_R[50], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_25 U1 (P[52], O_R[51], IN1_R[1], U__d1, U__d0, P[51]);
  U4DPPG_2_25 U2 (P[53], O_R[52], IN1_R[2], U__d1, U__d0, P[52]);
  U4DPPG_3_25 U3 (P[54], O_R[53], IN1_R[3], U__d1, U__d0, P[53]);
  U4DPPG_4_25 U4 (P[55], O_R[54], IN1_R[4], U__d1, U__d0, P[54]);
  U4DPPG_5_25 U5 (P[56], O_R[55], IN1_R[5], U__d1, U__d0, P[55]);
  U4DPPG_6_25 U6 (P[57], O_R[56], IN1_R[6], U__d1, U__d0, P[56]);
  U4DPPG_7_25 U7 (P[58], O_R[57], IN1_R[7], U__d1, U__d0, P[57]);
  U4DPPG_8_25 U8 (P[59], O_R[58], IN1_R[8], U__d1, U__d0, P[58]);
  U4DPPG_9_25 U9 (P[60], O_R[59], IN1_R[9], U__d1, U__d0, P[59]);
  U4DPPG_10_25 U10 (P[61], O_R[60], IN1_R[10], U__d1, U__d0, P[60]);
  U4DPPG_11_25 U11 (P[62], O_R[61], IN1_R[11], U__d1, U__d0, P[61]);
  U4DPPG_12_25 U12 (P[63], O_R[62], IN1_R[12], U__d1, U__d0, P[62]);
  U4DPPG_13_25 U13 (P[64], O_R[63], IN1_R[13], U__d1, U__d0, P[63]);
  U4DPPG_14_25 U14 (P[65], O_R[64], IN1_R[14], U__d1, U__d0, P[64]);
  U4DPPG_15_25 U15 (P[66], O_R[65], IN1_R[15], U__d1, U__d0, P[65]);
  U4DPPG_16_25 U16 (P[67], O_R[66], IN1_R[16], U__d1, U__d0, P[66]);
  U4DPPG_17_25 U17 (P[68], O_R[67], IN1_R[17], U__d1, U__d0, P[67]);
  U4DPPG_18_25 U18 (P[69], O_R[68], IN1_R[18], U__d1, U__d0, P[68]);
  U4DPPG_19_25 U19 (P[70], O_R[69], IN1_R[19], U__d1, U__d0, P[69]);
  U4DPPG_20_25 U20 (P[71], O_R[70], IN1_R[20], U__d1, U__d0, P[70]);
  U4DPPG_21_25 U21 (P[72], O_R[71], IN1_R[21], U__d1, U__d0, P[71]);
  U4DPPG_22_25 U22 (P[73], O_R[72], IN1_R[22], U__d1, U__d0, P[72]);
  U4DPPG_23_25 U23 (P[74], O_R[73], IN1_R[23], U__d1, U__d0, P[73]);
  U4DPPG_24_25 U24 (P[75], O_R[74], IN1_R[24], U__d1, U__d0, P[74]);
  U4DPPG_25_25 U25 (P[76], O_R[75], IN1_R[25], U__d1, U__d0, P[75]);
  U4DPPG_26_25 U26 (P[77], O_R[76], IN1_R[26], U__d1, U__d0, P[76]);
  U4DPPG_27_25 U27 (P[78], O_R[77], IN1_R[27], U__d1, U__d0, P[77]);
  U4DPPG_28_25 U28 (P[79], O_R[78], IN1_R[28], U__d1, U__d0, P[78]);
  U4DPPG_29_25 U29 (P[80], O_R[79], IN1_R[29], U__d1, U__d0, P[79]);
  U4DPPG_30_25 U30 (P[81], O_R[80], IN1_R[30], U__d1, U__d0, P[80]);
  U4DPPG_31_25 U31 (P[82], O_R[81], IN1_R[31], U__d1, U__d0, P[81]);
  U4DPPG_32_25 U32 (P[83], O_R[82], IN1_R[32], U__d1, U__d0, P[82]);
  U4DPPG_33_25 U33 (P[84], O_R[83], IN1_R[33], U__d1, U__d0, P[83]);
  U4DPPG_34_25 U34 (P[85], O_R[84], IN1_R[34], U__d1, U__d0, P[84]);
  U4DPPG_35_25 U35 (P[86], O_R[85], IN1_R[35], U__d1, U__d0, P[85]);
  U4DPPG_36_25 U36 (P[87], O_R[86], IN1_R[36], U__d1, U__d0, P[86]);
  U4DPPG_37_25 U37 (P[88], O_R[87], IN1_R[37], U__d1, U__d0, P[87]);
  U4DPPG_38_25 U38 (P[89], O_R[88], IN1_R[38], U__d1, U__d0, P[88]);
  U4DPPG_39_25 U39 (P[90], O_R[89], IN1_R[39], U__d1, U__d0, P[89]);
  U4DPPG_40_25 U40 (P[91], O_R[90], IN1_R[40], U__d1, U__d0, P[90]);
  U4DPPG_41_25 U41 (P[92], O_R[91], IN1_R[41], U__d1, U__d0, P[91]);
  U4DPPG_42_25 U42 (P[93], O_R[92], IN1_R[42], U__d1, U__d0, P[92]);
  U4DPPG_43_25 U43 (P[94], O_R[93], IN1_R[43], U__d1, U__d0, P[93]);
  U4DPPG_44_25 U44 (P[95], O_R[94], IN1_R[44], U__d1, U__d0, P[94]);
  U4DPPG_45_25 U45 (P[96], O_R[95], IN1_R[45], U__d1, U__d0, P[95]);
  U4DPPG_46_25 U46 (P[97], O_R[96], IN1_R[46], U__d1, U__d0, P[96]);
  U4DPPG_47_25 U47 (P[98], O_R[97], IN1_R[47], U__d1, U__d0, P[97]);
  U4DPPG_48_25 U48 (P[99], O_R[98], IN1_R[48], U__d1, U__d0, P[98]);
  U4DPPG_49_25 U49 (P[100], O_R[99], IN1_R[49], U__d1, U__d0, P[99]);
  U4DPPG_50_25 U50 (P[101], O_R[100], IN1_R[50], U__d1, U__d0, P[100]);
  U4DPPG_51_25 U51 (P[102], O_R[101], IN1_R[51], U__d1, U__d0, P[101]);
  U4DPPG_52_25 U52 (P[103], O_R[102], IN1_R[52], U__d1, U__d0, P[102]);
  U4DPPG_53_25 U53 (P[104], O_R[103], IN1_R[53], U__d1, U__d0, P[103]);
  U4DPPG_54_25 U54 (P[105], O_R[104], IN1_R[54], U__d1, U__d0, P[104]);
  U4DPPG_55_25 U55 (P[106], O_R[105], IN1_R[55], U__d1, U__d0, P[105]);
  U4DPPG_56_25 U56 (P[107], O_R[106], IN1_R[56], U__d1, U__d0, P[106]);
  U4DPPG_57_25 U57 (P[108], O_R[107], IN1_R[57], U__d1, U__d0, P[107]);
  U4DPPG_58_25 U58 (P[109], O_R[108], IN1_R[58], U__d1, U__d0, P[108]);
  U4DPPG_59_25 U59 (P[110], O_R[109], IN1_R[59], U__d1, U__d0, P[109]);
  U4DPPG_60_25 U60 (P[111], O_R[110], IN1_R[60], U__d1, U__d0, P[110]);
  U4DPPG_61_25 U61 (P[112], O_R[111], IN1_R[61], U__d1, U__d0, P[111]);
  U4DPPG_62_25 U62 (P[113], O_R[112], IN1_R[62], U__d1, U__d0, P[112]);
  U4DPPGH_63_25 U63 (O_T, O_R[113], IN1_T, U__d1, U__d0, P[113]);
endmodule

module TCU4VPPG_63_0_26 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [115:52] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [115:53] P;
  U4DPPGL_0_26 U0 (P[53], O_R[52], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_26 U1 (P[54], O_R[53], IN1_R[1], U__d1, U__d0, P[53]);
  U4DPPG_2_26 U2 (P[55], O_R[54], IN1_R[2], U__d1, U__d0, P[54]);
  U4DPPG_3_26 U3 (P[56], O_R[55], IN1_R[3], U__d1, U__d0, P[55]);
  U4DPPG_4_26 U4 (P[57], O_R[56], IN1_R[4], U__d1, U__d0, P[56]);
  U4DPPG_5_26 U5 (P[58], O_R[57], IN1_R[5], U__d1, U__d0, P[57]);
  U4DPPG_6_26 U6 (P[59], O_R[58], IN1_R[6], U__d1, U__d0, P[58]);
  U4DPPG_7_26 U7 (P[60], O_R[59], IN1_R[7], U__d1, U__d0, P[59]);
  U4DPPG_8_26 U8 (P[61], O_R[60], IN1_R[8], U__d1, U__d0, P[60]);
  U4DPPG_9_26 U9 (P[62], O_R[61], IN1_R[9], U__d1, U__d0, P[61]);
  U4DPPG_10_26 U10 (P[63], O_R[62], IN1_R[10], U__d1, U__d0, P[62]);
  U4DPPG_11_26 U11 (P[64], O_R[63], IN1_R[11], U__d1, U__d0, P[63]);
  U4DPPG_12_26 U12 (P[65], O_R[64], IN1_R[12], U__d1, U__d0, P[64]);
  U4DPPG_13_26 U13 (P[66], O_R[65], IN1_R[13], U__d1, U__d0, P[65]);
  U4DPPG_14_26 U14 (P[67], O_R[66], IN1_R[14], U__d1, U__d0, P[66]);
  U4DPPG_15_26 U15 (P[68], O_R[67], IN1_R[15], U__d1, U__d0, P[67]);
  U4DPPG_16_26 U16 (P[69], O_R[68], IN1_R[16], U__d1, U__d0, P[68]);
  U4DPPG_17_26 U17 (P[70], O_R[69], IN1_R[17], U__d1, U__d0, P[69]);
  U4DPPG_18_26 U18 (P[71], O_R[70], IN1_R[18], U__d1, U__d0, P[70]);
  U4DPPG_19_26 U19 (P[72], O_R[71], IN1_R[19], U__d1, U__d0, P[71]);
  U4DPPG_20_26 U20 (P[73], O_R[72], IN1_R[20], U__d1, U__d0, P[72]);
  U4DPPG_21_26 U21 (P[74], O_R[73], IN1_R[21], U__d1, U__d0, P[73]);
  U4DPPG_22_26 U22 (P[75], O_R[74], IN1_R[22], U__d1, U__d0, P[74]);
  U4DPPG_23_26 U23 (P[76], O_R[75], IN1_R[23], U__d1, U__d0, P[75]);
  U4DPPG_24_26 U24 (P[77], O_R[76], IN1_R[24], U__d1, U__d0, P[76]);
  U4DPPG_25_26 U25 (P[78], O_R[77], IN1_R[25], U__d1, U__d0, P[77]);
  U4DPPG_26_26 U26 (P[79], O_R[78], IN1_R[26], U__d1, U__d0, P[78]);
  U4DPPG_27_26 U27 (P[80], O_R[79], IN1_R[27], U__d1, U__d0, P[79]);
  U4DPPG_28_26 U28 (P[81], O_R[80], IN1_R[28], U__d1, U__d0, P[80]);
  U4DPPG_29_26 U29 (P[82], O_R[81], IN1_R[29], U__d1, U__d0, P[81]);
  U4DPPG_30_26 U30 (P[83], O_R[82], IN1_R[30], U__d1, U__d0, P[82]);
  U4DPPG_31_26 U31 (P[84], O_R[83], IN1_R[31], U__d1, U__d0, P[83]);
  U4DPPG_32_26 U32 (P[85], O_R[84], IN1_R[32], U__d1, U__d0, P[84]);
  U4DPPG_33_26 U33 (P[86], O_R[85], IN1_R[33], U__d1, U__d0, P[85]);
  U4DPPG_34_26 U34 (P[87], O_R[86], IN1_R[34], U__d1, U__d0, P[86]);
  U4DPPG_35_26 U35 (P[88], O_R[87], IN1_R[35], U__d1, U__d0, P[87]);
  U4DPPG_36_26 U36 (P[89], O_R[88], IN1_R[36], U__d1, U__d0, P[88]);
  U4DPPG_37_26 U37 (P[90], O_R[89], IN1_R[37], U__d1, U__d0, P[89]);
  U4DPPG_38_26 U38 (P[91], O_R[90], IN1_R[38], U__d1, U__d0, P[90]);
  U4DPPG_39_26 U39 (P[92], O_R[91], IN1_R[39], U__d1, U__d0, P[91]);
  U4DPPG_40_26 U40 (P[93], O_R[92], IN1_R[40], U__d1, U__d0, P[92]);
  U4DPPG_41_26 U41 (P[94], O_R[93], IN1_R[41], U__d1, U__d0, P[93]);
  U4DPPG_42_26 U42 (P[95], O_R[94], IN1_R[42], U__d1, U__d0, P[94]);
  U4DPPG_43_26 U43 (P[96], O_R[95], IN1_R[43], U__d1, U__d0, P[95]);
  U4DPPG_44_26 U44 (P[97], O_R[96], IN1_R[44], U__d1, U__d0, P[96]);
  U4DPPG_45_26 U45 (P[98], O_R[97], IN1_R[45], U__d1, U__d0, P[97]);
  U4DPPG_46_26 U46 (P[99], O_R[98], IN1_R[46], U__d1, U__d0, P[98]);
  U4DPPG_47_26 U47 (P[100], O_R[99], IN1_R[47], U__d1, U__d0, P[99]);
  U4DPPG_48_26 U48 (P[101], O_R[100], IN1_R[48], U__d1, U__d0, P[100]);
  U4DPPG_49_26 U49 (P[102], O_R[101], IN1_R[49], U__d1, U__d0, P[101]);
  U4DPPG_50_26 U50 (P[103], O_R[102], IN1_R[50], U__d1, U__d0, P[102]);
  U4DPPG_51_26 U51 (P[104], O_R[103], IN1_R[51], U__d1, U__d0, P[103]);
  U4DPPG_52_26 U52 (P[105], O_R[104], IN1_R[52], U__d1, U__d0, P[104]);
  U4DPPG_53_26 U53 (P[106], O_R[105], IN1_R[53], U__d1, U__d0, P[105]);
  U4DPPG_54_26 U54 (P[107], O_R[106], IN1_R[54], U__d1, U__d0, P[106]);
  U4DPPG_55_26 U55 (P[108], O_R[107], IN1_R[55], U__d1, U__d0, P[107]);
  U4DPPG_56_26 U56 (P[109], O_R[108], IN1_R[56], U__d1, U__d0, P[108]);
  U4DPPG_57_26 U57 (P[110], O_R[109], IN1_R[57], U__d1, U__d0, P[109]);
  U4DPPG_58_26 U58 (P[111], O_R[110], IN1_R[58], U__d1, U__d0, P[110]);
  U4DPPG_59_26 U59 (P[112], O_R[111], IN1_R[59], U__d1, U__d0, P[111]);
  U4DPPG_60_26 U60 (P[113], O_R[112], IN1_R[60], U__d1, U__d0, P[112]);
  U4DPPG_61_26 U61 (P[114], O_R[113], IN1_R[61], U__d1, U__d0, P[113]);
  U4DPPG_62_26 U62 (P[115], O_R[114], IN1_R[62], U__d1, U__d0, P[114]);
  U4DPPGH_63_26 U63 (O_T, O_R[115], IN1_T, U__d1, U__d0, P[115]);
endmodule

module TCU4VPPG_63_0_27 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [117:54] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [117:55] P;
  U4DPPGL_0_27 U0 (P[55], O_R[54], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_27 U1 (P[56], O_R[55], IN1_R[1], U__d1, U__d0, P[55]);
  U4DPPG_2_27 U2 (P[57], O_R[56], IN1_R[2], U__d1, U__d0, P[56]);
  U4DPPG_3_27 U3 (P[58], O_R[57], IN1_R[3], U__d1, U__d0, P[57]);
  U4DPPG_4_27 U4 (P[59], O_R[58], IN1_R[4], U__d1, U__d0, P[58]);
  U4DPPG_5_27 U5 (P[60], O_R[59], IN1_R[5], U__d1, U__d0, P[59]);
  U4DPPG_6_27 U6 (P[61], O_R[60], IN1_R[6], U__d1, U__d0, P[60]);
  U4DPPG_7_27 U7 (P[62], O_R[61], IN1_R[7], U__d1, U__d0, P[61]);
  U4DPPG_8_27 U8 (P[63], O_R[62], IN1_R[8], U__d1, U__d0, P[62]);
  U4DPPG_9_27 U9 (P[64], O_R[63], IN1_R[9], U__d1, U__d0, P[63]);
  U4DPPG_10_27 U10 (P[65], O_R[64], IN1_R[10], U__d1, U__d0, P[64]);
  U4DPPG_11_27 U11 (P[66], O_R[65], IN1_R[11], U__d1, U__d0, P[65]);
  U4DPPG_12_27 U12 (P[67], O_R[66], IN1_R[12], U__d1, U__d0, P[66]);
  U4DPPG_13_27 U13 (P[68], O_R[67], IN1_R[13], U__d1, U__d0, P[67]);
  U4DPPG_14_27 U14 (P[69], O_R[68], IN1_R[14], U__d1, U__d0, P[68]);
  U4DPPG_15_27 U15 (P[70], O_R[69], IN1_R[15], U__d1, U__d0, P[69]);
  U4DPPG_16_27 U16 (P[71], O_R[70], IN1_R[16], U__d1, U__d0, P[70]);
  U4DPPG_17_27 U17 (P[72], O_R[71], IN1_R[17], U__d1, U__d0, P[71]);
  U4DPPG_18_27 U18 (P[73], O_R[72], IN1_R[18], U__d1, U__d0, P[72]);
  U4DPPG_19_27 U19 (P[74], O_R[73], IN1_R[19], U__d1, U__d0, P[73]);
  U4DPPG_20_27 U20 (P[75], O_R[74], IN1_R[20], U__d1, U__d0, P[74]);
  U4DPPG_21_27 U21 (P[76], O_R[75], IN1_R[21], U__d1, U__d0, P[75]);
  U4DPPG_22_27 U22 (P[77], O_R[76], IN1_R[22], U__d1, U__d0, P[76]);
  U4DPPG_23_27 U23 (P[78], O_R[77], IN1_R[23], U__d1, U__d0, P[77]);
  U4DPPG_24_27 U24 (P[79], O_R[78], IN1_R[24], U__d1, U__d0, P[78]);
  U4DPPG_25_27 U25 (P[80], O_R[79], IN1_R[25], U__d1, U__d0, P[79]);
  U4DPPG_26_27 U26 (P[81], O_R[80], IN1_R[26], U__d1, U__d0, P[80]);
  U4DPPG_27_27 U27 (P[82], O_R[81], IN1_R[27], U__d1, U__d0, P[81]);
  U4DPPG_28_27 U28 (P[83], O_R[82], IN1_R[28], U__d1, U__d0, P[82]);
  U4DPPG_29_27 U29 (P[84], O_R[83], IN1_R[29], U__d1, U__d0, P[83]);
  U4DPPG_30_27 U30 (P[85], O_R[84], IN1_R[30], U__d1, U__d0, P[84]);
  U4DPPG_31_27 U31 (P[86], O_R[85], IN1_R[31], U__d1, U__d0, P[85]);
  U4DPPG_32_27 U32 (P[87], O_R[86], IN1_R[32], U__d1, U__d0, P[86]);
  U4DPPG_33_27 U33 (P[88], O_R[87], IN1_R[33], U__d1, U__d0, P[87]);
  U4DPPG_34_27 U34 (P[89], O_R[88], IN1_R[34], U__d1, U__d0, P[88]);
  U4DPPG_35_27 U35 (P[90], O_R[89], IN1_R[35], U__d1, U__d0, P[89]);
  U4DPPG_36_27 U36 (P[91], O_R[90], IN1_R[36], U__d1, U__d0, P[90]);
  U4DPPG_37_27 U37 (P[92], O_R[91], IN1_R[37], U__d1, U__d0, P[91]);
  U4DPPG_38_27 U38 (P[93], O_R[92], IN1_R[38], U__d1, U__d0, P[92]);
  U4DPPG_39_27 U39 (P[94], O_R[93], IN1_R[39], U__d1, U__d0, P[93]);
  U4DPPG_40_27 U40 (P[95], O_R[94], IN1_R[40], U__d1, U__d0, P[94]);
  U4DPPG_41_27 U41 (P[96], O_R[95], IN1_R[41], U__d1, U__d0, P[95]);
  U4DPPG_42_27 U42 (P[97], O_R[96], IN1_R[42], U__d1, U__d0, P[96]);
  U4DPPG_43_27 U43 (P[98], O_R[97], IN1_R[43], U__d1, U__d0, P[97]);
  U4DPPG_44_27 U44 (P[99], O_R[98], IN1_R[44], U__d1, U__d0, P[98]);
  U4DPPG_45_27 U45 (P[100], O_R[99], IN1_R[45], U__d1, U__d0, P[99]);
  U4DPPG_46_27 U46 (P[101], O_R[100], IN1_R[46], U__d1, U__d0, P[100]);
  U4DPPG_47_27 U47 (P[102], O_R[101], IN1_R[47], U__d1, U__d0, P[101]);
  U4DPPG_48_27 U48 (P[103], O_R[102], IN1_R[48], U__d1, U__d0, P[102]);
  U4DPPG_49_27 U49 (P[104], O_R[103], IN1_R[49], U__d1, U__d0, P[103]);
  U4DPPG_50_27 U50 (P[105], O_R[104], IN1_R[50], U__d1, U__d0, P[104]);
  U4DPPG_51_27 U51 (P[106], O_R[105], IN1_R[51], U__d1, U__d0, P[105]);
  U4DPPG_52_27 U52 (P[107], O_R[106], IN1_R[52], U__d1, U__d0, P[106]);
  U4DPPG_53_27 U53 (P[108], O_R[107], IN1_R[53], U__d1, U__d0, P[107]);
  U4DPPG_54_27 U54 (P[109], O_R[108], IN1_R[54], U__d1, U__d0, P[108]);
  U4DPPG_55_27 U55 (P[110], O_R[109], IN1_R[55], U__d1, U__d0, P[109]);
  U4DPPG_56_27 U56 (P[111], O_R[110], IN1_R[56], U__d1, U__d0, P[110]);
  U4DPPG_57_27 U57 (P[112], O_R[111], IN1_R[57], U__d1, U__d0, P[111]);
  U4DPPG_58_27 U58 (P[113], O_R[112], IN1_R[58], U__d1, U__d0, P[112]);
  U4DPPG_59_27 U59 (P[114], O_R[113], IN1_R[59], U__d1, U__d0, P[113]);
  U4DPPG_60_27 U60 (P[115], O_R[114], IN1_R[60], U__d1, U__d0, P[114]);
  U4DPPG_61_27 U61 (P[116], O_R[115], IN1_R[61], U__d1, U__d0, P[115]);
  U4DPPG_62_27 U62 (P[117], O_R[116], IN1_R[62], U__d1, U__d0, P[116]);
  U4DPPGH_63_27 U63 (O_T, O_R[117], IN1_T, U__d1, U__d0, P[117]);
endmodule

module TCU4VPPG_63_0_28 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [119:56] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [119:57] P;
  U4DPPGL_0_28 U0 (P[57], O_R[56], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_28 U1 (P[58], O_R[57], IN1_R[1], U__d1, U__d0, P[57]);
  U4DPPG_2_28 U2 (P[59], O_R[58], IN1_R[2], U__d1, U__d0, P[58]);
  U4DPPG_3_28 U3 (P[60], O_R[59], IN1_R[3], U__d1, U__d0, P[59]);
  U4DPPG_4_28 U4 (P[61], O_R[60], IN1_R[4], U__d1, U__d0, P[60]);
  U4DPPG_5_28 U5 (P[62], O_R[61], IN1_R[5], U__d1, U__d0, P[61]);
  U4DPPG_6_28 U6 (P[63], O_R[62], IN1_R[6], U__d1, U__d0, P[62]);
  U4DPPG_7_28 U7 (P[64], O_R[63], IN1_R[7], U__d1, U__d0, P[63]);
  U4DPPG_8_28 U8 (P[65], O_R[64], IN1_R[8], U__d1, U__d0, P[64]);
  U4DPPG_9_28 U9 (P[66], O_R[65], IN1_R[9], U__d1, U__d0, P[65]);
  U4DPPG_10_28 U10 (P[67], O_R[66], IN1_R[10], U__d1, U__d0, P[66]);
  U4DPPG_11_28 U11 (P[68], O_R[67], IN1_R[11], U__d1, U__d0, P[67]);
  U4DPPG_12_28 U12 (P[69], O_R[68], IN1_R[12], U__d1, U__d0, P[68]);
  U4DPPG_13_28 U13 (P[70], O_R[69], IN1_R[13], U__d1, U__d0, P[69]);
  U4DPPG_14_28 U14 (P[71], O_R[70], IN1_R[14], U__d1, U__d0, P[70]);
  U4DPPG_15_28 U15 (P[72], O_R[71], IN1_R[15], U__d1, U__d0, P[71]);
  U4DPPG_16_28 U16 (P[73], O_R[72], IN1_R[16], U__d1, U__d0, P[72]);
  U4DPPG_17_28 U17 (P[74], O_R[73], IN1_R[17], U__d1, U__d0, P[73]);
  U4DPPG_18_28 U18 (P[75], O_R[74], IN1_R[18], U__d1, U__d0, P[74]);
  U4DPPG_19_28 U19 (P[76], O_R[75], IN1_R[19], U__d1, U__d0, P[75]);
  U4DPPG_20_28 U20 (P[77], O_R[76], IN1_R[20], U__d1, U__d0, P[76]);
  U4DPPG_21_28 U21 (P[78], O_R[77], IN1_R[21], U__d1, U__d0, P[77]);
  U4DPPG_22_28 U22 (P[79], O_R[78], IN1_R[22], U__d1, U__d0, P[78]);
  U4DPPG_23_28 U23 (P[80], O_R[79], IN1_R[23], U__d1, U__d0, P[79]);
  U4DPPG_24_28 U24 (P[81], O_R[80], IN1_R[24], U__d1, U__d0, P[80]);
  U4DPPG_25_28 U25 (P[82], O_R[81], IN1_R[25], U__d1, U__d0, P[81]);
  U4DPPG_26_28 U26 (P[83], O_R[82], IN1_R[26], U__d1, U__d0, P[82]);
  U4DPPG_27_28 U27 (P[84], O_R[83], IN1_R[27], U__d1, U__d0, P[83]);
  U4DPPG_28_28 U28 (P[85], O_R[84], IN1_R[28], U__d1, U__d0, P[84]);
  U4DPPG_29_28 U29 (P[86], O_R[85], IN1_R[29], U__d1, U__d0, P[85]);
  U4DPPG_30_28 U30 (P[87], O_R[86], IN1_R[30], U__d1, U__d0, P[86]);
  U4DPPG_31_28 U31 (P[88], O_R[87], IN1_R[31], U__d1, U__d0, P[87]);
  U4DPPG_32_28 U32 (P[89], O_R[88], IN1_R[32], U__d1, U__d0, P[88]);
  U4DPPG_33_28 U33 (P[90], O_R[89], IN1_R[33], U__d1, U__d0, P[89]);
  U4DPPG_34_28 U34 (P[91], O_R[90], IN1_R[34], U__d1, U__d0, P[90]);
  U4DPPG_35_28 U35 (P[92], O_R[91], IN1_R[35], U__d1, U__d0, P[91]);
  U4DPPG_36_28 U36 (P[93], O_R[92], IN1_R[36], U__d1, U__d0, P[92]);
  U4DPPG_37_28 U37 (P[94], O_R[93], IN1_R[37], U__d1, U__d0, P[93]);
  U4DPPG_38_28 U38 (P[95], O_R[94], IN1_R[38], U__d1, U__d0, P[94]);
  U4DPPG_39_28 U39 (P[96], O_R[95], IN1_R[39], U__d1, U__d0, P[95]);
  U4DPPG_40_28 U40 (P[97], O_R[96], IN1_R[40], U__d1, U__d0, P[96]);
  U4DPPG_41_28 U41 (P[98], O_R[97], IN1_R[41], U__d1, U__d0, P[97]);
  U4DPPG_42_28 U42 (P[99], O_R[98], IN1_R[42], U__d1, U__d0, P[98]);
  U4DPPG_43_28 U43 (P[100], O_R[99], IN1_R[43], U__d1, U__d0, P[99]);
  U4DPPG_44_28 U44 (P[101], O_R[100], IN1_R[44], U__d1, U__d0, P[100]);
  U4DPPG_45_28 U45 (P[102], O_R[101], IN1_R[45], U__d1, U__d0, P[101]);
  U4DPPG_46_28 U46 (P[103], O_R[102], IN1_R[46], U__d1, U__d0, P[102]);
  U4DPPG_47_28 U47 (P[104], O_R[103], IN1_R[47], U__d1, U__d0, P[103]);
  U4DPPG_48_28 U48 (P[105], O_R[104], IN1_R[48], U__d1, U__d0, P[104]);
  U4DPPG_49_28 U49 (P[106], O_R[105], IN1_R[49], U__d1, U__d0, P[105]);
  U4DPPG_50_28 U50 (P[107], O_R[106], IN1_R[50], U__d1, U__d0, P[106]);
  U4DPPG_51_28 U51 (P[108], O_R[107], IN1_R[51], U__d1, U__d0, P[107]);
  U4DPPG_52_28 U52 (P[109], O_R[108], IN1_R[52], U__d1, U__d0, P[108]);
  U4DPPG_53_28 U53 (P[110], O_R[109], IN1_R[53], U__d1, U__d0, P[109]);
  U4DPPG_54_28 U54 (P[111], O_R[110], IN1_R[54], U__d1, U__d0, P[110]);
  U4DPPG_55_28 U55 (P[112], O_R[111], IN1_R[55], U__d1, U__d0, P[111]);
  U4DPPG_56_28 U56 (P[113], O_R[112], IN1_R[56], U__d1, U__d0, P[112]);
  U4DPPG_57_28 U57 (P[114], O_R[113], IN1_R[57], U__d1, U__d0, P[113]);
  U4DPPG_58_28 U58 (P[115], O_R[114], IN1_R[58], U__d1, U__d0, P[114]);
  U4DPPG_59_28 U59 (P[116], O_R[115], IN1_R[59], U__d1, U__d0, P[115]);
  U4DPPG_60_28 U60 (P[117], O_R[116], IN1_R[60], U__d1, U__d0, P[116]);
  U4DPPG_61_28 U61 (P[118], O_R[117], IN1_R[61], U__d1, U__d0, P[117]);
  U4DPPG_62_28 U62 (P[119], O_R[118], IN1_R[62], U__d1, U__d0, P[118]);
  U4DPPGH_63_28 U63 (O_T, O_R[119], IN1_T, U__d1, U__d0, P[119]);
endmodule

module TCU4VPPG_63_0_29 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [121:58] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [121:59] P;
  U4DPPGL_0_29 U0 (P[59], O_R[58], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_29 U1 (P[60], O_R[59], IN1_R[1], U__d1, U__d0, P[59]);
  U4DPPG_2_29 U2 (P[61], O_R[60], IN1_R[2], U__d1, U__d0, P[60]);
  U4DPPG_3_29 U3 (P[62], O_R[61], IN1_R[3], U__d1, U__d0, P[61]);
  U4DPPG_4_29 U4 (P[63], O_R[62], IN1_R[4], U__d1, U__d0, P[62]);
  U4DPPG_5_29 U5 (P[64], O_R[63], IN1_R[5], U__d1, U__d0, P[63]);
  U4DPPG_6_29 U6 (P[65], O_R[64], IN1_R[6], U__d1, U__d0, P[64]);
  U4DPPG_7_29 U7 (P[66], O_R[65], IN1_R[7], U__d1, U__d0, P[65]);
  U4DPPG_8_29 U8 (P[67], O_R[66], IN1_R[8], U__d1, U__d0, P[66]);
  U4DPPG_9_29 U9 (P[68], O_R[67], IN1_R[9], U__d1, U__d0, P[67]);
  U4DPPG_10_29 U10 (P[69], O_R[68], IN1_R[10], U__d1, U__d0, P[68]);
  U4DPPG_11_29 U11 (P[70], O_R[69], IN1_R[11], U__d1, U__d0, P[69]);
  U4DPPG_12_29 U12 (P[71], O_R[70], IN1_R[12], U__d1, U__d0, P[70]);
  U4DPPG_13_29 U13 (P[72], O_R[71], IN1_R[13], U__d1, U__d0, P[71]);
  U4DPPG_14_29 U14 (P[73], O_R[72], IN1_R[14], U__d1, U__d0, P[72]);
  U4DPPG_15_29 U15 (P[74], O_R[73], IN1_R[15], U__d1, U__d0, P[73]);
  U4DPPG_16_29 U16 (P[75], O_R[74], IN1_R[16], U__d1, U__d0, P[74]);
  U4DPPG_17_29 U17 (P[76], O_R[75], IN1_R[17], U__d1, U__d0, P[75]);
  U4DPPG_18_29 U18 (P[77], O_R[76], IN1_R[18], U__d1, U__d0, P[76]);
  U4DPPG_19_29 U19 (P[78], O_R[77], IN1_R[19], U__d1, U__d0, P[77]);
  U4DPPG_20_29 U20 (P[79], O_R[78], IN1_R[20], U__d1, U__d0, P[78]);
  U4DPPG_21_29 U21 (P[80], O_R[79], IN1_R[21], U__d1, U__d0, P[79]);
  U4DPPG_22_29 U22 (P[81], O_R[80], IN1_R[22], U__d1, U__d0, P[80]);
  U4DPPG_23_29 U23 (P[82], O_R[81], IN1_R[23], U__d1, U__d0, P[81]);
  U4DPPG_24_29 U24 (P[83], O_R[82], IN1_R[24], U__d1, U__d0, P[82]);
  U4DPPG_25_29 U25 (P[84], O_R[83], IN1_R[25], U__d1, U__d0, P[83]);
  U4DPPG_26_29 U26 (P[85], O_R[84], IN1_R[26], U__d1, U__d0, P[84]);
  U4DPPG_27_29 U27 (P[86], O_R[85], IN1_R[27], U__d1, U__d0, P[85]);
  U4DPPG_28_29 U28 (P[87], O_R[86], IN1_R[28], U__d1, U__d0, P[86]);
  U4DPPG_29_29 U29 (P[88], O_R[87], IN1_R[29], U__d1, U__d0, P[87]);
  U4DPPG_30_29 U30 (P[89], O_R[88], IN1_R[30], U__d1, U__d0, P[88]);
  U4DPPG_31_29 U31 (P[90], O_R[89], IN1_R[31], U__d1, U__d0, P[89]);
  U4DPPG_32_29 U32 (P[91], O_R[90], IN1_R[32], U__d1, U__d0, P[90]);
  U4DPPG_33_29 U33 (P[92], O_R[91], IN1_R[33], U__d1, U__d0, P[91]);
  U4DPPG_34_29 U34 (P[93], O_R[92], IN1_R[34], U__d1, U__d0, P[92]);
  U4DPPG_35_29 U35 (P[94], O_R[93], IN1_R[35], U__d1, U__d0, P[93]);
  U4DPPG_36_29 U36 (P[95], O_R[94], IN1_R[36], U__d1, U__d0, P[94]);
  U4DPPG_37_29 U37 (P[96], O_R[95], IN1_R[37], U__d1, U__d0, P[95]);
  U4DPPG_38_29 U38 (P[97], O_R[96], IN1_R[38], U__d1, U__d0, P[96]);
  U4DPPG_39_29 U39 (P[98], O_R[97], IN1_R[39], U__d1, U__d0, P[97]);
  U4DPPG_40_29 U40 (P[99], O_R[98], IN1_R[40], U__d1, U__d0, P[98]);
  U4DPPG_41_29 U41 (P[100], O_R[99], IN1_R[41], U__d1, U__d0, P[99]);
  U4DPPG_42_29 U42 (P[101], O_R[100], IN1_R[42], U__d1, U__d0, P[100]);
  U4DPPG_43_29 U43 (P[102], O_R[101], IN1_R[43], U__d1, U__d0, P[101]);
  U4DPPG_44_29 U44 (P[103], O_R[102], IN1_R[44], U__d1, U__d0, P[102]);
  U4DPPG_45_29 U45 (P[104], O_R[103], IN1_R[45], U__d1, U__d0, P[103]);
  U4DPPG_46_29 U46 (P[105], O_R[104], IN1_R[46], U__d1, U__d0, P[104]);
  U4DPPG_47_29 U47 (P[106], O_R[105], IN1_R[47], U__d1, U__d0, P[105]);
  U4DPPG_48_29 U48 (P[107], O_R[106], IN1_R[48], U__d1, U__d0, P[106]);
  U4DPPG_49_29 U49 (P[108], O_R[107], IN1_R[49], U__d1, U__d0, P[107]);
  U4DPPG_50_29 U50 (P[109], O_R[108], IN1_R[50], U__d1, U__d0, P[108]);
  U4DPPG_51_29 U51 (P[110], O_R[109], IN1_R[51], U__d1, U__d0, P[109]);
  U4DPPG_52_29 U52 (P[111], O_R[110], IN1_R[52], U__d1, U__d0, P[110]);
  U4DPPG_53_29 U53 (P[112], O_R[111], IN1_R[53], U__d1, U__d0, P[111]);
  U4DPPG_54_29 U54 (P[113], O_R[112], IN1_R[54], U__d1, U__d0, P[112]);
  U4DPPG_55_29 U55 (P[114], O_R[113], IN1_R[55], U__d1, U__d0, P[113]);
  U4DPPG_56_29 U56 (P[115], O_R[114], IN1_R[56], U__d1, U__d0, P[114]);
  U4DPPG_57_29 U57 (P[116], O_R[115], IN1_R[57], U__d1, U__d0, P[115]);
  U4DPPG_58_29 U58 (P[117], O_R[116], IN1_R[58], U__d1, U__d0, P[116]);
  U4DPPG_59_29 U59 (P[118], O_R[117], IN1_R[59], U__d1, U__d0, P[117]);
  U4DPPG_60_29 U60 (P[119], O_R[118], IN1_R[60], U__d1, U__d0, P[118]);
  U4DPPG_61_29 U61 (P[120], O_R[119], IN1_R[61], U__d1, U__d0, P[119]);
  U4DPPG_62_29 U62 (P[121], O_R[120], IN1_R[62], U__d1, U__d0, P[120]);
  U4DPPGH_63_29 U63 (O_T, O_R[121], IN1_T, U__d1, U__d0, P[121]);
endmodule

module TCU4VPPG_63_0_3 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [69:6] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [69:7] P;
  U4DPPGL_0_3 U0 (P[7], O_R[6], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_3 U1 (P[8], O_R[7], IN1_R[1], U__d1, U__d0, P[7]);
  U4DPPG_2_3 U2 (P[9], O_R[8], IN1_R[2], U__d1, U__d0, P[8]);
  U4DPPG_3_3 U3 (P[10], O_R[9], IN1_R[3], U__d1, U__d0, P[9]);
  U4DPPG_4_3 U4 (P[11], O_R[10], IN1_R[4], U__d1, U__d0, P[10]);
  U4DPPG_5_3 U5 (P[12], O_R[11], IN1_R[5], U__d1, U__d0, P[11]);
  U4DPPG_6_3 U6 (P[13], O_R[12], IN1_R[6], U__d1, U__d0, P[12]);
  U4DPPG_7_3 U7 (P[14], O_R[13], IN1_R[7], U__d1, U__d0, P[13]);
  U4DPPG_8_3 U8 (P[15], O_R[14], IN1_R[8], U__d1, U__d0, P[14]);
  U4DPPG_9_3 U9 (P[16], O_R[15], IN1_R[9], U__d1, U__d0, P[15]);
  U4DPPG_10_3 U10 (P[17], O_R[16], IN1_R[10], U__d1, U__d0, P[16]);
  U4DPPG_11_3 U11 (P[18], O_R[17], IN1_R[11], U__d1, U__d0, P[17]);
  U4DPPG_12_3 U12 (P[19], O_R[18], IN1_R[12], U__d1, U__d0, P[18]);
  U4DPPG_13_3 U13 (P[20], O_R[19], IN1_R[13], U__d1, U__d0, P[19]);
  U4DPPG_14_3 U14 (P[21], O_R[20], IN1_R[14], U__d1, U__d0, P[20]);
  U4DPPG_15_3 U15 (P[22], O_R[21], IN1_R[15], U__d1, U__d0, P[21]);
  U4DPPG_16_3 U16 (P[23], O_R[22], IN1_R[16], U__d1, U__d0, P[22]);
  U4DPPG_17_3 U17 (P[24], O_R[23], IN1_R[17], U__d1, U__d0, P[23]);
  U4DPPG_18_3 U18 (P[25], O_R[24], IN1_R[18], U__d1, U__d0, P[24]);
  U4DPPG_19_3 U19 (P[26], O_R[25], IN1_R[19], U__d1, U__d0, P[25]);
  U4DPPG_20_3 U20 (P[27], O_R[26], IN1_R[20], U__d1, U__d0, P[26]);
  U4DPPG_21_3 U21 (P[28], O_R[27], IN1_R[21], U__d1, U__d0, P[27]);
  U4DPPG_22_3 U22 (P[29], O_R[28], IN1_R[22], U__d1, U__d0, P[28]);
  U4DPPG_23_3 U23 (P[30], O_R[29], IN1_R[23], U__d1, U__d0, P[29]);
  U4DPPG_24_3 U24 (P[31], O_R[30], IN1_R[24], U__d1, U__d0, P[30]);
  U4DPPG_25_3 U25 (P[32], O_R[31], IN1_R[25], U__d1, U__d0, P[31]);
  U4DPPG_26_3 U26 (P[33], O_R[32], IN1_R[26], U__d1, U__d0, P[32]);
  U4DPPG_27_3 U27 (P[34], O_R[33], IN1_R[27], U__d1, U__d0, P[33]);
  U4DPPG_28_3 U28 (P[35], O_R[34], IN1_R[28], U__d1, U__d0, P[34]);
  U4DPPG_29_3 U29 (P[36], O_R[35], IN1_R[29], U__d1, U__d0, P[35]);
  U4DPPG_30_3 U30 (P[37], O_R[36], IN1_R[30], U__d1, U__d0, P[36]);
  U4DPPG_31_3 U31 (P[38], O_R[37], IN1_R[31], U__d1, U__d0, P[37]);
  U4DPPG_32_3 U32 (P[39], O_R[38], IN1_R[32], U__d1, U__d0, P[38]);
  U4DPPG_33_3 U33 (P[40], O_R[39], IN1_R[33], U__d1, U__d0, P[39]);
  U4DPPG_34_3 U34 (P[41], O_R[40], IN1_R[34], U__d1, U__d0, P[40]);
  U4DPPG_35_3 U35 (P[42], O_R[41], IN1_R[35], U__d1, U__d0, P[41]);
  U4DPPG_36_3 U36 (P[43], O_R[42], IN1_R[36], U__d1, U__d0, P[42]);
  U4DPPG_37_3 U37 (P[44], O_R[43], IN1_R[37], U__d1, U__d0, P[43]);
  U4DPPG_38_3 U38 (P[45], O_R[44], IN1_R[38], U__d1, U__d0, P[44]);
  U4DPPG_39_3 U39 (P[46], O_R[45], IN1_R[39], U__d1, U__d0, P[45]);
  U4DPPG_40_3 U40 (P[47], O_R[46], IN1_R[40], U__d1, U__d0, P[46]);
  U4DPPG_41_3 U41 (P[48], O_R[47], IN1_R[41], U__d1, U__d0, P[47]);
  U4DPPG_42_3 U42 (P[49], O_R[48], IN1_R[42], U__d1, U__d0, P[48]);
  U4DPPG_43_3 U43 (P[50], O_R[49], IN1_R[43], U__d1, U__d0, P[49]);
  U4DPPG_44_3 U44 (P[51], O_R[50], IN1_R[44], U__d1, U__d0, P[50]);
  U4DPPG_45_3 U45 (P[52], O_R[51], IN1_R[45], U__d1, U__d0, P[51]);
  U4DPPG_46_3 U46 (P[53], O_R[52], IN1_R[46], U__d1, U__d0, P[52]);
  U4DPPG_47_3 U47 (P[54], O_R[53], IN1_R[47], U__d1, U__d0, P[53]);
  U4DPPG_48_3 U48 (P[55], O_R[54], IN1_R[48], U__d1, U__d0, P[54]);
  U4DPPG_49_3 U49 (P[56], O_R[55], IN1_R[49], U__d1, U__d0, P[55]);
  U4DPPG_50_3 U50 (P[57], O_R[56], IN1_R[50], U__d1, U__d0, P[56]);
  U4DPPG_51_3 U51 (P[58], O_R[57], IN1_R[51], U__d1, U__d0, P[57]);
  U4DPPG_52_3 U52 (P[59], O_R[58], IN1_R[52], U__d1, U__d0, P[58]);
  U4DPPG_53_3 U53 (P[60], O_R[59], IN1_R[53], U__d1, U__d0, P[59]);
  U4DPPG_54_3 U54 (P[61], O_R[60], IN1_R[54], U__d1, U__d0, P[60]);
  U4DPPG_55_3 U55 (P[62], O_R[61], IN1_R[55], U__d1, U__d0, P[61]);
  U4DPPG_56_3 U56 (P[63], O_R[62], IN1_R[56], U__d1, U__d0, P[62]);
  U4DPPG_57_3 U57 (P[64], O_R[63], IN1_R[57], U__d1, U__d0, P[63]);
  U4DPPG_58_3 U58 (P[65], O_R[64], IN1_R[58], U__d1, U__d0, P[64]);
  U4DPPG_59_3 U59 (P[66], O_R[65], IN1_R[59], U__d1, U__d0, P[65]);
  U4DPPG_60_3 U60 (P[67], O_R[66], IN1_R[60], U__d1, U__d0, P[66]);
  U4DPPG_61_3 U61 (P[68], O_R[67], IN1_R[61], U__d1, U__d0, P[67]);
  U4DPPG_62_3 U62 (P[69], O_R[68], IN1_R[62], U__d1, U__d0, P[68]);
  U4DPPGH_63_3 U63 (O_T, O_R[69], IN1_T, U__d1, U__d0, P[69]);
endmodule

module TCU4VPPG_63_0_30 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [123:60] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [123:61] P;
  U4DPPGL_0_30 U0 (P[61], O_R[60], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_30 U1 (P[62], O_R[61], IN1_R[1], U__d1, U__d0, P[61]);
  U4DPPG_2_30 U2 (P[63], O_R[62], IN1_R[2], U__d1, U__d0, P[62]);
  U4DPPG_3_30 U3 (P[64], O_R[63], IN1_R[3], U__d1, U__d0, P[63]);
  U4DPPG_4_30 U4 (P[65], O_R[64], IN1_R[4], U__d1, U__d0, P[64]);
  U4DPPG_5_30 U5 (P[66], O_R[65], IN1_R[5], U__d1, U__d0, P[65]);
  U4DPPG_6_30 U6 (P[67], O_R[66], IN1_R[6], U__d1, U__d0, P[66]);
  U4DPPG_7_30 U7 (P[68], O_R[67], IN1_R[7], U__d1, U__d0, P[67]);
  U4DPPG_8_30 U8 (P[69], O_R[68], IN1_R[8], U__d1, U__d0, P[68]);
  U4DPPG_9_30 U9 (P[70], O_R[69], IN1_R[9], U__d1, U__d0, P[69]);
  U4DPPG_10_30 U10 (P[71], O_R[70], IN1_R[10], U__d1, U__d0, P[70]);
  U4DPPG_11_30 U11 (P[72], O_R[71], IN1_R[11], U__d1, U__d0, P[71]);
  U4DPPG_12_30 U12 (P[73], O_R[72], IN1_R[12], U__d1, U__d0, P[72]);
  U4DPPG_13_30 U13 (P[74], O_R[73], IN1_R[13], U__d1, U__d0, P[73]);
  U4DPPG_14_30 U14 (P[75], O_R[74], IN1_R[14], U__d1, U__d0, P[74]);
  U4DPPG_15_30 U15 (P[76], O_R[75], IN1_R[15], U__d1, U__d0, P[75]);
  U4DPPG_16_30 U16 (P[77], O_R[76], IN1_R[16], U__d1, U__d0, P[76]);
  U4DPPG_17_30 U17 (P[78], O_R[77], IN1_R[17], U__d1, U__d0, P[77]);
  U4DPPG_18_30 U18 (P[79], O_R[78], IN1_R[18], U__d1, U__d0, P[78]);
  U4DPPG_19_30 U19 (P[80], O_R[79], IN1_R[19], U__d1, U__d0, P[79]);
  U4DPPG_20_30 U20 (P[81], O_R[80], IN1_R[20], U__d1, U__d0, P[80]);
  U4DPPG_21_30 U21 (P[82], O_R[81], IN1_R[21], U__d1, U__d0, P[81]);
  U4DPPG_22_30 U22 (P[83], O_R[82], IN1_R[22], U__d1, U__d0, P[82]);
  U4DPPG_23_30 U23 (P[84], O_R[83], IN1_R[23], U__d1, U__d0, P[83]);
  U4DPPG_24_30 U24 (P[85], O_R[84], IN1_R[24], U__d1, U__d0, P[84]);
  U4DPPG_25_30 U25 (P[86], O_R[85], IN1_R[25], U__d1, U__d0, P[85]);
  U4DPPG_26_30 U26 (P[87], O_R[86], IN1_R[26], U__d1, U__d0, P[86]);
  U4DPPG_27_30 U27 (P[88], O_R[87], IN1_R[27], U__d1, U__d0, P[87]);
  U4DPPG_28_30 U28 (P[89], O_R[88], IN1_R[28], U__d1, U__d0, P[88]);
  U4DPPG_29_30 U29 (P[90], O_R[89], IN1_R[29], U__d1, U__d0, P[89]);
  U4DPPG_30_30 U30 (P[91], O_R[90], IN1_R[30], U__d1, U__d0, P[90]);
  U4DPPG_31_30 U31 (P[92], O_R[91], IN1_R[31], U__d1, U__d0, P[91]);
  U4DPPG_32_30 U32 (P[93], O_R[92], IN1_R[32], U__d1, U__d0, P[92]);
  U4DPPG_33_30 U33 (P[94], O_R[93], IN1_R[33], U__d1, U__d0, P[93]);
  U4DPPG_34_30 U34 (P[95], O_R[94], IN1_R[34], U__d1, U__d0, P[94]);
  U4DPPG_35_30 U35 (P[96], O_R[95], IN1_R[35], U__d1, U__d0, P[95]);
  U4DPPG_36_30 U36 (P[97], O_R[96], IN1_R[36], U__d1, U__d0, P[96]);
  U4DPPG_37_30 U37 (P[98], O_R[97], IN1_R[37], U__d1, U__d0, P[97]);
  U4DPPG_38_30 U38 (P[99], O_R[98], IN1_R[38], U__d1, U__d0, P[98]);
  U4DPPG_39_30 U39 (P[100], O_R[99], IN1_R[39], U__d1, U__d0, P[99]);
  U4DPPG_40_30 U40 (P[101], O_R[100], IN1_R[40], U__d1, U__d0, P[100]);
  U4DPPG_41_30 U41 (P[102], O_R[101], IN1_R[41], U__d1, U__d0, P[101]);
  U4DPPG_42_30 U42 (P[103], O_R[102], IN1_R[42], U__d1, U__d0, P[102]);
  U4DPPG_43_30 U43 (P[104], O_R[103], IN1_R[43], U__d1, U__d0, P[103]);
  U4DPPG_44_30 U44 (P[105], O_R[104], IN1_R[44], U__d1, U__d0, P[104]);
  U4DPPG_45_30 U45 (P[106], O_R[105], IN1_R[45], U__d1, U__d0, P[105]);
  U4DPPG_46_30 U46 (P[107], O_R[106], IN1_R[46], U__d1, U__d0, P[106]);
  U4DPPG_47_30 U47 (P[108], O_R[107], IN1_R[47], U__d1, U__d0, P[107]);
  U4DPPG_48_30 U48 (P[109], O_R[108], IN1_R[48], U__d1, U__d0, P[108]);
  U4DPPG_49_30 U49 (P[110], O_R[109], IN1_R[49], U__d1, U__d0, P[109]);
  U4DPPG_50_30 U50 (P[111], O_R[110], IN1_R[50], U__d1, U__d0, P[110]);
  U4DPPG_51_30 U51 (P[112], O_R[111], IN1_R[51], U__d1, U__d0, P[111]);
  U4DPPG_52_30 U52 (P[113], O_R[112], IN1_R[52], U__d1, U__d0, P[112]);
  U4DPPG_53_30 U53 (P[114], O_R[113], IN1_R[53], U__d1, U__d0, P[113]);
  U4DPPG_54_30 U54 (P[115], O_R[114], IN1_R[54], U__d1, U__d0, P[114]);
  U4DPPG_55_30 U55 (P[116], O_R[115], IN1_R[55], U__d1, U__d0, P[115]);
  U4DPPG_56_30 U56 (P[117], O_R[116], IN1_R[56], U__d1, U__d0, P[116]);
  U4DPPG_57_30 U57 (P[118], O_R[117], IN1_R[57], U__d1, U__d0, P[117]);
  U4DPPG_58_30 U58 (P[119], O_R[118], IN1_R[58], U__d1, U__d0, P[118]);
  U4DPPG_59_30 U59 (P[120], O_R[119], IN1_R[59], U__d1, U__d0, P[119]);
  U4DPPG_60_30 U60 (P[121], O_R[120], IN1_R[60], U__d1, U__d0, P[120]);
  U4DPPG_61_30 U61 (P[122], O_R[121], IN1_R[61], U__d1, U__d0, P[121]);
  U4DPPG_62_30 U62 (P[123], O_R[122], IN1_R[62], U__d1, U__d0, P[122]);
  U4DPPGH_63_30 U63 (O_T, O_R[123], IN1_T, U__d1, U__d0, P[123]);
endmodule

module TCU4VPPG_63_0_31 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [125:62] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [125:63] P;
  U4DPPGL_0_31 U0 (P[63], O_R[62], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_31 U1 (P[64], O_R[63], IN1_R[1], U__d1, U__d0, P[63]);
  U4DPPG_2_31 U2 (P[65], O_R[64], IN1_R[2], U__d1, U__d0, P[64]);
  U4DPPG_3_31 U3 (P[66], O_R[65], IN1_R[3], U__d1, U__d0, P[65]);
  U4DPPG_4_31 U4 (P[67], O_R[66], IN1_R[4], U__d1, U__d0, P[66]);
  U4DPPG_5_31 U5 (P[68], O_R[67], IN1_R[5], U__d1, U__d0, P[67]);
  U4DPPG_6_31 U6 (P[69], O_R[68], IN1_R[6], U__d1, U__d0, P[68]);
  U4DPPG_7_31 U7 (P[70], O_R[69], IN1_R[7], U__d1, U__d0, P[69]);
  U4DPPG_8_31 U8 (P[71], O_R[70], IN1_R[8], U__d1, U__d0, P[70]);
  U4DPPG_9_31 U9 (P[72], O_R[71], IN1_R[9], U__d1, U__d0, P[71]);
  U4DPPG_10_31 U10 (P[73], O_R[72], IN1_R[10], U__d1, U__d0, P[72]);
  U4DPPG_11_31 U11 (P[74], O_R[73], IN1_R[11], U__d1, U__d0, P[73]);
  U4DPPG_12_31 U12 (P[75], O_R[74], IN1_R[12], U__d1, U__d0, P[74]);
  U4DPPG_13_31 U13 (P[76], O_R[75], IN1_R[13], U__d1, U__d0, P[75]);
  U4DPPG_14_31 U14 (P[77], O_R[76], IN1_R[14], U__d1, U__d0, P[76]);
  U4DPPG_15_31 U15 (P[78], O_R[77], IN1_R[15], U__d1, U__d0, P[77]);
  U4DPPG_16_31 U16 (P[79], O_R[78], IN1_R[16], U__d1, U__d0, P[78]);
  U4DPPG_17_31 U17 (P[80], O_R[79], IN1_R[17], U__d1, U__d0, P[79]);
  U4DPPG_18_31 U18 (P[81], O_R[80], IN1_R[18], U__d1, U__d0, P[80]);
  U4DPPG_19_31 U19 (P[82], O_R[81], IN1_R[19], U__d1, U__d0, P[81]);
  U4DPPG_20_31 U20 (P[83], O_R[82], IN1_R[20], U__d1, U__d0, P[82]);
  U4DPPG_21_31 U21 (P[84], O_R[83], IN1_R[21], U__d1, U__d0, P[83]);
  U4DPPG_22_31 U22 (P[85], O_R[84], IN1_R[22], U__d1, U__d0, P[84]);
  U4DPPG_23_31 U23 (P[86], O_R[85], IN1_R[23], U__d1, U__d0, P[85]);
  U4DPPG_24_31 U24 (P[87], O_R[86], IN1_R[24], U__d1, U__d0, P[86]);
  U4DPPG_25_31 U25 (P[88], O_R[87], IN1_R[25], U__d1, U__d0, P[87]);
  U4DPPG_26_31 U26 (P[89], O_R[88], IN1_R[26], U__d1, U__d0, P[88]);
  U4DPPG_27_31 U27 (P[90], O_R[89], IN1_R[27], U__d1, U__d0, P[89]);
  U4DPPG_28_31 U28 (P[91], O_R[90], IN1_R[28], U__d1, U__d0, P[90]);
  U4DPPG_29_31 U29 (P[92], O_R[91], IN1_R[29], U__d1, U__d0, P[91]);
  U4DPPG_30_31 U30 (P[93], O_R[92], IN1_R[30], U__d1, U__d0, P[92]);
  U4DPPG_31_31 U31 (P[94], O_R[93], IN1_R[31], U__d1, U__d0, P[93]);
  U4DPPG_32_31 U32 (P[95], O_R[94], IN1_R[32], U__d1, U__d0, P[94]);
  U4DPPG_33_31 U33 (P[96], O_R[95], IN1_R[33], U__d1, U__d0, P[95]);
  U4DPPG_34_31 U34 (P[97], O_R[96], IN1_R[34], U__d1, U__d0, P[96]);
  U4DPPG_35_31 U35 (P[98], O_R[97], IN1_R[35], U__d1, U__d0, P[97]);
  U4DPPG_36_31 U36 (P[99], O_R[98], IN1_R[36], U__d1, U__d0, P[98]);
  U4DPPG_37_31 U37 (P[100], O_R[99], IN1_R[37], U__d1, U__d0, P[99]);
  U4DPPG_38_31 U38 (P[101], O_R[100], IN1_R[38], U__d1, U__d0, P[100]);
  U4DPPG_39_31 U39 (P[102], O_R[101], IN1_R[39], U__d1, U__d0, P[101]);
  U4DPPG_40_31 U40 (P[103], O_R[102], IN1_R[40], U__d1, U__d0, P[102]);
  U4DPPG_41_31 U41 (P[104], O_R[103], IN1_R[41], U__d1, U__d0, P[103]);
  U4DPPG_42_31 U42 (P[105], O_R[104], IN1_R[42], U__d1, U__d0, P[104]);
  U4DPPG_43_31 U43 (P[106], O_R[105], IN1_R[43], U__d1, U__d0, P[105]);
  U4DPPG_44_31 U44 (P[107], O_R[106], IN1_R[44], U__d1, U__d0, P[106]);
  U4DPPG_45_31 U45 (P[108], O_R[107], IN1_R[45], U__d1, U__d0, P[107]);
  U4DPPG_46_31 U46 (P[109], O_R[108], IN1_R[46], U__d1, U__d0, P[108]);
  U4DPPG_47_31 U47 (P[110], O_R[109], IN1_R[47], U__d1, U__d0, P[109]);
  U4DPPG_48_31 U48 (P[111], O_R[110], IN1_R[48], U__d1, U__d0, P[110]);
  U4DPPG_49_31 U49 (P[112], O_R[111], IN1_R[49], U__d1, U__d0, P[111]);
  U4DPPG_50_31 U50 (P[113], O_R[112], IN1_R[50], U__d1, U__d0, P[112]);
  U4DPPG_51_31 U51 (P[114], O_R[113], IN1_R[51], U__d1, U__d0, P[113]);
  U4DPPG_52_31 U52 (P[115], O_R[114], IN1_R[52], U__d1, U__d0, P[114]);
  U4DPPG_53_31 U53 (P[116], O_R[115], IN1_R[53], U__d1, U__d0, P[115]);
  U4DPPG_54_31 U54 (P[117], O_R[116], IN1_R[54], U__d1, U__d0, P[116]);
  U4DPPG_55_31 U55 (P[118], O_R[117], IN1_R[55], U__d1, U__d0, P[117]);
  U4DPPG_56_31 U56 (P[119], O_R[118], IN1_R[56], U__d1, U__d0, P[118]);
  U4DPPG_57_31 U57 (P[120], O_R[119], IN1_R[57], U__d1, U__d0, P[119]);
  U4DPPG_58_31 U58 (P[121], O_R[120], IN1_R[58], U__d1, U__d0, P[120]);
  U4DPPG_59_31 U59 (P[122], O_R[121], IN1_R[59], U__d1, U__d0, P[121]);
  U4DPPG_60_31 U60 (P[123], O_R[122], IN1_R[60], U__d1, U__d0, P[122]);
  U4DPPG_61_31 U61 (P[124], O_R[123], IN1_R[61], U__d1, U__d0, P[123]);
  U4DPPG_62_31 U62 (P[125], O_R[124], IN1_R[62], U__d1, U__d0, P[124]);
  U4DPPGH_63_31 U63 (O_T, O_R[125], IN1_T, U__d1, U__d0, P[125]);
endmodule

module TCU4VPPG_63_0_4 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [71:8] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [71:9] P;
  U4DPPGL_0_4 U0 (P[9], O_R[8], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_4 U1 (P[10], O_R[9], IN1_R[1], U__d1, U__d0, P[9]);
  U4DPPG_2_4 U2 (P[11], O_R[10], IN1_R[2], U__d1, U__d0, P[10]);
  U4DPPG_3_4 U3 (P[12], O_R[11], IN1_R[3], U__d1, U__d0, P[11]);
  U4DPPG_4_4 U4 (P[13], O_R[12], IN1_R[4], U__d1, U__d0, P[12]);
  U4DPPG_5_4 U5 (P[14], O_R[13], IN1_R[5], U__d1, U__d0, P[13]);
  U4DPPG_6_4 U6 (P[15], O_R[14], IN1_R[6], U__d1, U__d0, P[14]);
  U4DPPG_7_4 U7 (P[16], O_R[15], IN1_R[7], U__d1, U__d0, P[15]);
  U4DPPG_8_4 U8 (P[17], O_R[16], IN1_R[8], U__d1, U__d0, P[16]);
  U4DPPG_9_4 U9 (P[18], O_R[17], IN1_R[9], U__d1, U__d0, P[17]);
  U4DPPG_10_4 U10 (P[19], O_R[18], IN1_R[10], U__d1, U__d0, P[18]);
  U4DPPG_11_4 U11 (P[20], O_R[19], IN1_R[11], U__d1, U__d0, P[19]);
  U4DPPG_12_4 U12 (P[21], O_R[20], IN1_R[12], U__d1, U__d0, P[20]);
  U4DPPG_13_4 U13 (P[22], O_R[21], IN1_R[13], U__d1, U__d0, P[21]);
  U4DPPG_14_4 U14 (P[23], O_R[22], IN1_R[14], U__d1, U__d0, P[22]);
  U4DPPG_15_4 U15 (P[24], O_R[23], IN1_R[15], U__d1, U__d0, P[23]);
  U4DPPG_16_4 U16 (P[25], O_R[24], IN1_R[16], U__d1, U__d0, P[24]);
  U4DPPG_17_4 U17 (P[26], O_R[25], IN1_R[17], U__d1, U__d0, P[25]);
  U4DPPG_18_4 U18 (P[27], O_R[26], IN1_R[18], U__d1, U__d0, P[26]);
  U4DPPG_19_4 U19 (P[28], O_R[27], IN1_R[19], U__d1, U__d0, P[27]);
  U4DPPG_20_4 U20 (P[29], O_R[28], IN1_R[20], U__d1, U__d0, P[28]);
  U4DPPG_21_4 U21 (P[30], O_R[29], IN1_R[21], U__d1, U__d0, P[29]);
  U4DPPG_22_4 U22 (P[31], O_R[30], IN1_R[22], U__d1, U__d0, P[30]);
  U4DPPG_23_4 U23 (P[32], O_R[31], IN1_R[23], U__d1, U__d0, P[31]);
  U4DPPG_24_4 U24 (P[33], O_R[32], IN1_R[24], U__d1, U__d0, P[32]);
  U4DPPG_25_4 U25 (P[34], O_R[33], IN1_R[25], U__d1, U__d0, P[33]);
  U4DPPG_26_4 U26 (P[35], O_R[34], IN1_R[26], U__d1, U__d0, P[34]);
  U4DPPG_27_4 U27 (P[36], O_R[35], IN1_R[27], U__d1, U__d0, P[35]);
  U4DPPG_28_4 U28 (P[37], O_R[36], IN1_R[28], U__d1, U__d0, P[36]);
  U4DPPG_29_4 U29 (P[38], O_R[37], IN1_R[29], U__d1, U__d0, P[37]);
  U4DPPG_30_4 U30 (P[39], O_R[38], IN1_R[30], U__d1, U__d0, P[38]);
  U4DPPG_31_4 U31 (P[40], O_R[39], IN1_R[31], U__d1, U__d0, P[39]);
  U4DPPG_32_4 U32 (P[41], O_R[40], IN1_R[32], U__d1, U__d0, P[40]);
  U4DPPG_33_4 U33 (P[42], O_R[41], IN1_R[33], U__d1, U__d0, P[41]);
  U4DPPG_34_4 U34 (P[43], O_R[42], IN1_R[34], U__d1, U__d0, P[42]);
  U4DPPG_35_4 U35 (P[44], O_R[43], IN1_R[35], U__d1, U__d0, P[43]);
  U4DPPG_36_4 U36 (P[45], O_R[44], IN1_R[36], U__d1, U__d0, P[44]);
  U4DPPG_37_4 U37 (P[46], O_R[45], IN1_R[37], U__d1, U__d0, P[45]);
  U4DPPG_38_4 U38 (P[47], O_R[46], IN1_R[38], U__d1, U__d0, P[46]);
  U4DPPG_39_4 U39 (P[48], O_R[47], IN1_R[39], U__d1, U__d0, P[47]);
  U4DPPG_40_4 U40 (P[49], O_R[48], IN1_R[40], U__d1, U__d0, P[48]);
  U4DPPG_41_4 U41 (P[50], O_R[49], IN1_R[41], U__d1, U__d0, P[49]);
  U4DPPG_42_4 U42 (P[51], O_R[50], IN1_R[42], U__d1, U__d0, P[50]);
  U4DPPG_43_4 U43 (P[52], O_R[51], IN1_R[43], U__d1, U__d0, P[51]);
  U4DPPG_44_4 U44 (P[53], O_R[52], IN1_R[44], U__d1, U__d0, P[52]);
  U4DPPG_45_4 U45 (P[54], O_R[53], IN1_R[45], U__d1, U__d0, P[53]);
  U4DPPG_46_4 U46 (P[55], O_R[54], IN1_R[46], U__d1, U__d0, P[54]);
  U4DPPG_47_4 U47 (P[56], O_R[55], IN1_R[47], U__d1, U__d0, P[55]);
  U4DPPG_48_4 U48 (P[57], O_R[56], IN1_R[48], U__d1, U__d0, P[56]);
  U4DPPG_49_4 U49 (P[58], O_R[57], IN1_R[49], U__d1, U__d0, P[57]);
  U4DPPG_50_4 U50 (P[59], O_R[58], IN1_R[50], U__d1, U__d0, P[58]);
  U4DPPG_51_4 U51 (P[60], O_R[59], IN1_R[51], U__d1, U__d0, P[59]);
  U4DPPG_52_4 U52 (P[61], O_R[60], IN1_R[52], U__d1, U__d0, P[60]);
  U4DPPG_53_4 U53 (P[62], O_R[61], IN1_R[53], U__d1, U__d0, P[61]);
  U4DPPG_54_4 U54 (P[63], O_R[62], IN1_R[54], U__d1, U__d0, P[62]);
  U4DPPG_55_4 U55 (P[64], O_R[63], IN1_R[55], U__d1, U__d0, P[63]);
  U4DPPG_56_4 U56 (P[65], O_R[64], IN1_R[56], U__d1, U__d0, P[64]);
  U4DPPG_57_4 U57 (P[66], O_R[65], IN1_R[57], U__d1, U__d0, P[65]);
  U4DPPG_58_4 U58 (P[67], O_R[66], IN1_R[58], U__d1, U__d0, P[66]);
  U4DPPG_59_4 U59 (P[68], O_R[67], IN1_R[59], U__d1, U__d0, P[67]);
  U4DPPG_60_4 U60 (P[69], O_R[68], IN1_R[60], U__d1, U__d0, P[68]);
  U4DPPG_61_4 U61 (P[70], O_R[69], IN1_R[61], U__d1, U__d0, P[69]);
  U4DPPG_62_4 U62 (P[71], O_R[70], IN1_R[62], U__d1, U__d0, P[70]);
  U4DPPGH_63_4 U63 (O_T, O_R[71], IN1_T, U__d1, U__d0, P[71]);
endmodule

module TCU4VPPG_63_0_5 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [73:10] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [73:11] P;
  U4DPPGL_0_5 U0 (P[11], O_R[10], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_5 U1 (P[12], O_R[11], IN1_R[1], U__d1, U__d0, P[11]);
  U4DPPG_2_5 U2 (P[13], O_R[12], IN1_R[2], U__d1, U__d0, P[12]);
  U4DPPG_3_5 U3 (P[14], O_R[13], IN1_R[3], U__d1, U__d0, P[13]);
  U4DPPG_4_5 U4 (P[15], O_R[14], IN1_R[4], U__d1, U__d0, P[14]);
  U4DPPG_5_5 U5 (P[16], O_R[15], IN1_R[5], U__d1, U__d0, P[15]);
  U4DPPG_6_5 U6 (P[17], O_R[16], IN1_R[6], U__d1, U__d0, P[16]);
  U4DPPG_7_5 U7 (P[18], O_R[17], IN1_R[7], U__d1, U__d0, P[17]);
  U4DPPG_8_5 U8 (P[19], O_R[18], IN1_R[8], U__d1, U__d0, P[18]);
  U4DPPG_9_5 U9 (P[20], O_R[19], IN1_R[9], U__d1, U__d0, P[19]);
  U4DPPG_10_5 U10 (P[21], O_R[20], IN1_R[10], U__d1, U__d0, P[20]);
  U4DPPG_11_5 U11 (P[22], O_R[21], IN1_R[11], U__d1, U__d0, P[21]);
  U4DPPG_12_5 U12 (P[23], O_R[22], IN1_R[12], U__d1, U__d0, P[22]);
  U4DPPG_13_5 U13 (P[24], O_R[23], IN1_R[13], U__d1, U__d0, P[23]);
  U4DPPG_14_5 U14 (P[25], O_R[24], IN1_R[14], U__d1, U__d0, P[24]);
  U4DPPG_15_5 U15 (P[26], O_R[25], IN1_R[15], U__d1, U__d0, P[25]);
  U4DPPG_16_5 U16 (P[27], O_R[26], IN1_R[16], U__d1, U__d0, P[26]);
  U4DPPG_17_5 U17 (P[28], O_R[27], IN1_R[17], U__d1, U__d0, P[27]);
  U4DPPG_18_5 U18 (P[29], O_R[28], IN1_R[18], U__d1, U__d0, P[28]);
  U4DPPG_19_5 U19 (P[30], O_R[29], IN1_R[19], U__d1, U__d0, P[29]);
  U4DPPG_20_5 U20 (P[31], O_R[30], IN1_R[20], U__d1, U__d0, P[30]);
  U4DPPG_21_5 U21 (P[32], O_R[31], IN1_R[21], U__d1, U__d0, P[31]);
  U4DPPG_22_5 U22 (P[33], O_R[32], IN1_R[22], U__d1, U__d0, P[32]);
  U4DPPG_23_5 U23 (P[34], O_R[33], IN1_R[23], U__d1, U__d0, P[33]);
  U4DPPG_24_5 U24 (P[35], O_R[34], IN1_R[24], U__d1, U__d0, P[34]);
  U4DPPG_25_5 U25 (P[36], O_R[35], IN1_R[25], U__d1, U__d0, P[35]);
  U4DPPG_26_5 U26 (P[37], O_R[36], IN1_R[26], U__d1, U__d0, P[36]);
  U4DPPG_27_5 U27 (P[38], O_R[37], IN1_R[27], U__d1, U__d0, P[37]);
  U4DPPG_28_5 U28 (P[39], O_R[38], IN1_R[28], U__d1, U__d0, P[38]);
  U4DPPG_29_5 U29 (P[40], O_R[39], IN1_R[29], U__d1, U__d0, P[39]);
  U4DPPG_30_5 U30 (P[41], O_R[40], IN1_R[30], U__d1, U__d0, P[40]);
  U4DPPG_31_5 U31 (P[42], O_R[41], IN1_R[31], U__d1, U__d0, P[41]);
  U4DPPG_32_5 U32 (P[43], O_R[42], IN1_R[32], U__d1, U__d0, P[42]);
  U4DPPG_33_5 U33 (P[44], O_R[43], IN1_R[33], U__d1, U__d0, P[43]);
  U4DPPG_34_5 U34 (P[45], O_R[44], IN1_R[34], U__d1, U__d0, P[44]);
  U4DPPG_35_5 U35 (P[46], O_R[45], IN1_R[35], U__d1, U__d0, P[45]);
  U4DPPG_36_5 U36 (P[47], O_R[46], IN1_R[36], U__d1, U__d0, P[46]);
  U4DPPG_37_5 U37 (P[48], O_R[47], IN1_R[37], U__d1, U__d0, P[47]);
  U4DPPG_38_5 U38 (P[49], O_R[48], IN1_R[38], U__d1, U__d0, P[48]);
  U4DPPG_39_5 U39 (P[50], O_R[49], IN1_R[39], U__d1, U__d0, P[49]);
  U4DPPG_40_5 U40 (P[51], O_R[50], IN1_R[40], U__d1, U__d0, P[50]);
  U4DPPG_41_5 U41 (P[52], O_R[51], IN1_R[41], U__d1, U__d0, P[51]);
  U4DPPG_42_5 U42 (P[53], O_R[52], IN1_R[42], U__d1, U__d0, P[52]);
  U4DPPG_43_5 U43 (P[54], O_R[53], IN1_R[43], U__d1, U__d0, P[53]);
  U4DPPG_44_5 U44 (P[55], O_R[54], IN1_R[44], U__d1, U__d0, P[54]);
  U4DPPG_45_5 U45 (P[56], O_R[55], IN1_R[45], U__d1, U__d0, P[55]);
  U4DPPG_46_5 U46 (P[57], O_R[56], IN1_R[46], U__d1, U__d0, P[56]);
  U4DPPG_47_5 U47 (P[58], O_R[57], IN1_R[47], U__d1, U__d0, P[57]);
  U4DPPG_48_5 U48 (P[59], O_R[58], IN1_R[48], U__d1, U__d0, P[58]);
  U4DPPG_49_5 U49 (P[60], O_R[59], IN1_R[49], U__d1, U__d0, P[59]);
  U4DPPG_50_5 U50 (P[61], O_R[60], IN1_R[50], U__d1, U__d0, P[60]);
  U4DPPG_51_5 U51 (P[62], O_R[61], IN1_R[51], U__d1, U__d0, P[61]);
  U4DPPG_52_5 U52 (P[63], O_R[62], IN1_R[52], U__d1, U__d0, P[62]);
  U4DPPG_53_5 U53 (P[64], O_R[63], IN1_R[53], U__d1, U__d0, P[63]);
  U4DPPG_54_5 U54 (P[65], O_R[64], IN1_R[54], U__d1, U__d0, P[64]);
  U4DPPG_55_5 U55 (P[66], O_R[65], IN1_R[55], U__d1, U__d0, P[65]);
  U4DPPG_56_5 U56 (P[67], O_R[66], IN1_R[56], U__d1, U__d0, P[66]);
  U4DPPG_57_5 U57 (P[68], O_R[67], IN1_R[57], U__d1, U__d0, P[67]);
  U4DPPG_58_5 U58 (P[69], O_R[68], IN1_R[58], U__d1, U__d0, P[68]);
  U4DPPG_59_5 U59 (P[70], O_R[69], IN1_R[59], U__d1, U__d0, P[69]);
  U4DPPG_60_5 U60 (P[71], O_R[70], IN1_R[60], U__d1, U__d0, P[70]);
  U4DPPG_61_5 U61 (P[72], O_R[71], IN1_R[61], U__d1, U__d0, P[71]);
  U4DPPG_62_5 U62 (P[73], O_R[72], IN1_R[62], U__d1, U__d0, P[72]);
  U4DPPGH_63_5 U63 (O_T, O_R[73], IN1_T, U__d1, U__d0, P[73]);
endmodule

module TCU4VPPG_63_0_6 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [75:12] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [75:13] P;
  U4DPPGL_0_6 U0 (P[13], O_R[12], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_6 U1 (P[14], O_R[13], IN1_R[1], U__d1, U__d0, P[13]);
  U4DPPG_2_6 U2 (P[15], O_R[14], IN1_R[2], U__d1, U__d0, P[14]);
  U4DPPG_3_6 U3 (P[16], O_R[15], IN1_R[3], U__d1, U__d0, P[15]);
  U4DPPG_4_6 U4 (P[17], O_R[16], IN1_R[4], U__d1, U__d0, P[16]);
  U4DPPG_5_6 U5 (P[18], O_R[17], IN1_R[5], U__d1, U__d0, P[17]);
  U4DPPG_6_6 U6 (P[19], O_R[18], IN1_R[6], U__d1, U__d0, P[18]);
  U4DPPG_7_6 U7 (P[20], O_R[19], IN1_R[7], U__d1, U__d0, P[19]);
  U4DPPG_8_6 U8 (P[21], O_R[20], IN1_R[8], U__d1, U__d0, P[20]);
  U4DPPG_9_6 U9 (P[22], O_R[21], IN1_R[9], U__d1, U__d0, P[21]);
  U4DPPG_10_6 U10 (P[23], O_R[22], IN1_R[10], U__d1, U__d0, P[22]);
  U4DPPG_11_6 U11 (P[24], O_R[23], IN1_R[11], U__d1, U__d0, P[23]);
  U4DPPG_12_6 U12 (P[25], O_R[24], IN1_R[12], U__d1, U__d0, P[24]);
  U4DPPG_13_6 U13 (P[26], O_R[25], IN1_R[13], U__d1, U__d0, P[25]);
  U4DPPG_14_6 U14 (P[27], O_R[26], IN1_R[14], U__d1, U__d0, P[26]);
  U4DPPG_15_6 U15 (P[28], O_R[27], IN1_R[15], U__d1, U__d0, P[27]);
  U4DPPG_16_6 U16 (P[29], O_R[28], IN1_R[16], U__d1, U__d0, P[28]);
  U4DPPG_17_6 U17 (P[30], O_R[29], IN1_R[17], U__d1, U__d0, P[29]);
  U4DPPG_18_6 U18 (P[31], O_R[30], IN1_R[18], U__d1, U__d0, P[30]);
  U4DPPG_19_6 U19 (P[32], O_R[31], IN1_R[19], U__d1, U__d0, P[31]);
  U4DPPG_20_6 U20 (P[33], O_R[32], IN1_R[20], U__d1, U__d0, P[32]);
  U4DPPG_21_6 U21 (P[34], O_R[33], IN1_R[21], U__d1, U__d0, P[33]);
  U4DPPG_22_6 U22 (P[35], O_R[34], IN1_R[22], U__d1, U__d0, P[34]);
  U4DPPG_23_6 U23 (P[36], O_R[35], IN1_R[23], U__d1, U__d0, P[35]);
  U4DPPG_24_6 U24 (P[37], O_R[36], IN1_R[24], U__d1, U__d0, P[36]);
  U4DPPG_25_6 U25 (P[38], O_R[37], IN1_R[25], U__d1, U__d0, P[37]);
  U4DPPG_26_6 U26 (P[39], O_R[38], IN1_R[26], U__d1, U__d0, P[38]);
  U4DPPG_27_6 U27 (P[40], O_R[39], IN1_R[27], U__d1, U__d0, P[39]);
  U4DPPG_28_6 U28 (P[41], O_R[40], IN1_R[28], U__d1, U__d0, P[40]);
  U4DPPG_29_6 U29 (P[42], O_R[41], IN1_R[29], U__d1, U__d0, P[41]);
  U4DPPG_30_6 U30 (P[43], O_R[42], IN1_R[30], U__d1, U__d0, P[42]);
  U4DPPG_31_6 U31 (P[44], O_R[43], IN1_R[31], U__d1, U__d0, P[43]);
  U4DPPG_32_6 U32 (P[45], O_R[44], IN1_R[32], U__d1, U__d0, P[44]);
  U4DPPG_33_6 U33 (P[46], O_R[45], IN1_R[33], U__d1, U__d0, P[45]);
  U4DPPG_34_6 U34 (P[47], O_R[46], IN1_R[34], U__d1, U__d0, P[46]);
  U4DPPG_35_6 U35 (P[48], O_R[47], IN1_R[35], U__d1, U__d0, P[47]);
  U4DPPG_36_6 U36 (P[49], O_R[48], IN1_R[36], U__d1, U__d0, P[48]);
  U4DPPG_37_6 U37 (P[50], O_R[49], IN1_R[37], U__d1, U__d0, P[49]);
  U4DPPG_38_6 U38 (P[51], O_R[50], IN1_R[38], U__d1, U__d0, P[50]);
  U4DPPG_39_6 U39 (P[52], O_R[51], IN1_R[39], U__d1, U__d0, P[51]);
  U4DPPG_40_6 U40 (P[53], O_R[52], IN1_R[40], U__d1, U__d0, P[52]);
  U4DPPG_41_6 U41 (P[54], O_R[53], IN1_R[41], U__d1, U__d0, P[53]);
  U4DPPG_42_6 U42 (P[55], O_R[54], IN1_R[42], U__d1, U__d0, P[54]);
  U4DPPG_43_6 U43 (P[56], O_R[55], IN1_R[43], U__d1, U__d0, P[55]);
  U4DPPG_44_6 U44 (P[57], O_R[56], IN1_R[44], U__d1, U__d0, P[56]);
  U4DPPG_45_6 U45 (P[58], O_R[57], IN1_R[45], U__d1, U__d0, P[57]);
  U4DPPG_46_6 U46 (P[59], O_R[58], IN1_R[46], U__d1, U__d0, P[58]);
  U4DPPG_47_6 U47 (P[60], O_R[59], IN1_R[47], U__d1, U__d0, P[59]);
  U4DPPG_48_6 U48 (P[61], O_R[60], IN1_R[48], U__d1, U__d0, P[60]);
  U4DPPG_49_6 U49 (P[62], O_R[61], IN1_R[49], U__d1, U__d0, P[61]);
  U4DPPG_50_6 U50 (P[63], O_R[62], IN1_R[50], U__d1, U__d0, P[62]);
  U4DPPG_51_6 U51 (P[64], O_R[63], IN1_R[51], U__d1, U__d0, P[63]);
  U4DPPG_52_6 U52 (P[65], O_R[64], IN1_R[52], U__d1, U__d0, P[64]);
  U4DPPG_53_6 U53 (P[66], O_R[65], IN1_R[53], U__d1, U__d0, P[65]);
  U4DPPG_54_6 U54 (P[67], O_R[66], IN1_R[54], U__d1, U__d0, P[66]);
  U4DPPG_55_6 U55 (P[68], O_R[67], IN1_R[55], U__d1, U__d0, P[67]);
  U4DPPG_56_6 U56 (P[69], O_R[68], IN1_R[56], U__d1, U__d0, P[68]);
  U4DPPG_57_6 U57 (P[70], O_R[69], IN1_R[57], U__d1, U__d0, P[69]);
  U4DPPG_58_6 U58 (P[71], O_R[70], IN1_R[58], U__d1, U__d0, P[70]);
  U4DPPG_59_6 U59 (P[72], O_R[71], IN1_R[59], U__d1, U__d0, P[71]);
  U4DPPG_60_6 U60 (P[73], O_R[72], IN1_R[60], U__d1, U__d0, P[72]);
  U4DPPG_61_6 U61 (P[74], O_R[73], IN1_R[61], U__d1, U__d0, P[73]);
  U4DPPG_62_6 U62 (P[75], O_R[74], IN1_R[62], U__d1, U__d0, P[74]);
  U4DPPGH_63_6 U63 (O_T, O_R[75], IN1_T, U__d1, U__d0, P[75]);
endmodule

module TCU4VPPG_63_0_7 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [77:14] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [77:15] P;
  U4DPPGL_0_7 U0 (P[15], O_R[14], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_7 U1 (P[16], O_R[15], IN1_R[1], U__d1, U__d0, P[15]);
  U4DPPG_2_7 U2 (P[17], O_R[16], IN1_R[2], U__d1, U__d0, P[16]);
  U4DPPG_3_7 U3 (P[18], O_R[17], IN1_R[3], U__d1, U__d0, P[17]);
  U4DPPG_4_7 U4 (P[19], O_R[18], IN1_R[4], U__d1, U__d0, P[18]);
  U4DPPG_5_7 U5 (P[20], O_R[19], IN1_R[5], U__d1, U__d0, P[19]);
  U4DPPG_6_7 U6 (P[21], O_R[20], IN1_R[6], U__d1, U__d0, P[20]);
  U4DPPG_7_7 U7 (P[22], O_R[21], IN1_R[7], U__d1, U__d0, P[21]);
  U4DPPG_8_7 U8 (P[23], O_R[22], IN1_R[8], U__d1, U__d0, P[22]);
  U4DPPG_9_7 U9 (P[24], O_R[23], IN1_R[9], U__d1, U__d0, P[23]);
  U4DPPG_10_7 U10 (P[25], O_R[24], IN1_R[10], U__d1, U__d0, P[24]);
  U4DPPG_11_7 U11 (P[26], O_R[25], IN1_R[11], U__d1, U__d0, P[25]);
  U4DPPG_12_7 U12 (P[27], O_R[26], IN1_R[12], U__d1, U__d0, P[26]);
  U4DPPG_13_7 U13 (P[28], O_R[27], IN1_R[13], U__d1, U__d0, P[27]);
  U4DPPG_14_7 U14 (P[29], O_R[28], IN1_R[14], U__d1, U__d0, P[28]);
  U4DPPG_15_7 U15 (P[30], O_R[29], IN1_R[15], U__d1, U__d0, P[29]);
  U4DPPG_16_7 U16 (P[31], O_R[30], IN1_R[16], U__d1, U__d0, P[30]);
  U4DPPG_17_7 U17 (P[32], O_R[31], IN1_R[17], U__d1, U__d0, P[31]);
  U4DPPG_18_7 U18 (P[33], O_R[32], IN1_R[18], U__d1, U__d0, P[32]);
  U4DPPG_19_7 U19 (P[34], O_R[33], IN1_R[19], U__d1, U__d0, P[33]);
  U4DPPG_20_7 U20 (P[35], O_R[34], IN1_R[20], U__d1, U__d0, P[34]);
  U4DPPG_21_7 U21 (P[36], O_R[35], IN1_R[21], U__d1, U__d0, P[35]);
  U4DPPG_22_7 U22 (P[37], O_R[36], IN1_R[22], U__d1, U__d0, P[36]);
  U4DPPG_23_7 U23 (P[38], O_R[37], IN1_R[23], U__d1, U__d0, P[37]);
  U4DPPG_24_7 U24 (P[39], O_R[38], IN1_R[24], U__d1, U__d0, P[38]);
  U4DPPG_25_7 U25 (P[40], O_R[39], IN1_R[25], U__d1, U__d0, P[39]);
  U4DPPG_26_7 U26 (P[41], O_R[40], IN1_R[26], U__d1, U__d0, P[40]);
  U4DPPG_27_7 U27 (P[42], O_R[41], IN1_R[27], U__d1, U__d0, P[41]);
  U4DPPG_28_7 U28 (P[43], O_R[42], IN1_R[28], U__d1, U__d0, P[42]);
  U4DPPG_29_7 U29 (P[44], O_R[43], IN1_R[29], U__d1, U__d0, P[43]);
  U4DPPG_30_7 U30 (P[45], O_R[44], IN1_R[30], U__d1, U__d0, P[44]);
  U4DPPG_31_7 U31 (P[46], O_R[45], IN1_R[31], U__d1, U__d0, P[45]);
  U4DPPG_32_7 U32 (P[47], O_R[46], IN1_R[32], U__d1, U__d0, P[46]);
  U4DPPG_33_7 U33 (P[48], O_R[47], IN1_R[33], U__d1, U__d0, P[47]);
  U4DPPG_34_7 U34 (P[49], O_R[48], IN1_R[34], U__d1, U__d0, P[48]);
  U4DPPG_35_7 U35 (P[50], O_R[49], IN1_R[35], U__d1, U__d0, P[49]);
  U4DPPG_36_7 U36 (P[51], O_R[50], IN1_R[36], U__d1, U__d0, P[50]);
  U4DPPG_37_7 U37 (P[52], O_R[51], IN1_R[37], U__d1, U__d0, P[51]);
  U4DPPG_38_7 U38 (P[53], O_R[52], IN1_R[38], U__d1, U__d0, P[52]);
  U4DPPG_39_7 U39 (P[54], O_R[53], IN1_R[39], U__d1, U__d0, P[53]);
  U4DPPG_40_7 U40 (P[55], O_R[54], IN1_R[40], U__d1, U__d0, P[54]);
  U4DPPG_41_7 U41 (P[56], O_R[55], IN1_R[41], U__d1, U__d0, P[55]);
  U4DPPG_42_7 U42 (P[57], O_R[56], IN1_R[42], U__d1, U__d0, P[56]);
  U4DPPG_43_7 U43 (P[58], O_R[57], IN1_R[43], U__d1, U__d0, P[57]);
  U4DPPG_44_7 U44 (P[59], O_R[58], IN1_R[44], U__d1, U__d0, P[58]);
  U4DPPG_45_7 U45 (P[60], O_R[59], IN1_R[45], U__d1, U__d0, P[59]);
  U4DPPG_46_7 U46 (P[61], O_R[60], IN1_R[46], U__d1, U__d0, P[60]);
  U4DPPG_47_7 U47 (P[62], O_R[61], IN1_R[47], U__d1, U__d0, P[61]);
  U4DPPG_48_7 U48 (P[63], O_R[62], IN1_R[48], U__d1, U__d0, P[62]);
  U4DPPG_49_7 U49 (P[64], O_R[63], IN1_R[49], U__d1, U__d0, P[63]);
  U4DPPG_50_7 U50 (P[65], O_R[64], IN1_R[50], U__d1, U__d0, P[64]);
  U4DPPG_51_7 U51 (P[66], O_R[65], IN1_R[51], U__d1, U__d0, P[65]);
  U4DPPG_52_7 U52 (P[67], O_R[66], IN1_R[52], U__d1, U__d0, P[66]);
  U4DPPG_53_7 U53 (P[68], O_R[67], IN1_R[53], U__d1, U__d0, P[67]);
  U4DPPG_54_7 U54 (P[69], O_R[68], IN1_R[54], U__d1, U__d0, P[68]);
  U4DPPG_55_7 U55 (P[70], O_R[69], IN1_R[55], U__d1, U__d0, P[69]);
  U4DPPG_56_7 U56 (P[71], O_R[70], IN1_R[56], U__d1, U__d0, P[70]);
  U4DPPG_57_7 U57 (P[72], O_R[71], IN1_R[57], U__d1, U__d0, P[71]);
  U4DPPG_58_7 U58 (P[73], O_R[72], IN1_R[58], U__d1, U__d0, P[72]);
  U4DPPG_59_7 U59 (P[74], O_R[73], IN1_R[59], U__d1, U__d0, P[73]);
  U4DPPG_60_7 U60 (P[75], O_R[74], IN1_R[60], U__d1, U__d0, P[74]);
  U4DPPG_61_7 U61 (P[76], O_R[75], IN1_R[61], U__d1, U__d0, P[75]);
  U4DPPG_62_7 U62 (P[77], O_R[76], IN1_R[62], U__d1, U__d0, P[76]);
  U4DPPGH_63_7 U63 (O_T, O_R[77], IN1_T, U__d1, U__d0, P[77]);
endmodule

module TCU4VPPG_63_0_8 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [79:16] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [79:17] P;
  U4DPPGL_0_8 U0 (P[17], O_R[16], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_8 U1 (P[18], O_R[17], IN1_R[1], U__d1, U__d0, P[17]);
  U4DPPG_2_8 U2 (P[19], O_R[18], IN1_R[2], U__d1, U__d0, P[18]);
  U4DPPG_3_8 U3 (P[20], O_R[19], IN1_R[3], U__d1, U__d0, P[19]);
  U4DPPG_4_8 U4 (P[21], O_R[20], IN1_R[4], U__d1, U__d0, P[20]);
  U4DPPG_5_8 U5 (P[22], O_R[21], IN1_R[5], U__d1, U__d0, P[21]);
  U4DPPG_6_8 U6 (P[23], O_R[22], IN1_R[6], U__d1, U__d0, P[22]);
  U4DPPG_7_8 U7 (P[24], O_R[23], IN1_R[7], U__d1, U__d0, P[23]);
  U4DPPG_8_8 U8 (P[25], O_R[24], IN1_R[8], U__d1, U__d0, P[24]);
  U4DPPG_9_8 U9 (P[26], O_R[25], IN1_R[9], U__d1, U__d0, P[25]);
  U4DPPG_10_8 U10 (P[27], O_R[26], IN1_R[10], U__d1, U__d0, P[26]);
  U4DPPG_11_8 U11 (P[28], O_R[27], IN1_R[11], U__d1, U__d0, P[27]);
  U4DPPG_12_8 U12 (P[29], O_R[28], IN1_R[12], U__d1, U__d0, P[28]);
  U4DPPG_13_8 U13 (P[30], O_R[29], IN1_R[13], U__d1, U__d0, P[29]);
  U4DPPG_14_8 U14 (P[31], O_R[30], IN1_R[14], U__d1, U__d0, P[30]);
  U4DPPG_15_8 U15 (P[32], O_R[31], IN1_R[15], U__d1, U__d0, P[31]);
  U4DPPG_16_8 U16 (P[33], O_R[32], IN1_R[16], U__d1, U__d0, P[32]);
  U4DPPG_17_8 U17 (P[34], O_R[33], IN1_R[17], U__d1, U__d0, P[33]);
  U4DPPG_18_8 U18 (P[35], O_R[34], IN1_R[18], U__d1, U__d0, P[34]);
  U4DPPG_19_8 U19 (P[36], O_R[35], IN1_R[19], U__d1, U__d0, P[35]);
  U4DPPG_20_8 U20 (P[37], O_R[36], IN1_R[20], U__d1, U__d0, P[36]);
  U4DPPG_21_8 U21 (P[38], O_R[37], IN1_R[21], U__d1, U__d0, P[37]);
  U4DPPG_22_8 U22 (P[39], O_R[38], IN1_R[22], U__d1, U__d0, P[38]);
  U4DPPG_23_8 U23 (P[40], O_R[39], IN1_R[23], U__d1, U__d0, P[39]);
  U4DPPG_24_8 U24 (P[41], O_R[40], IN1_R[24], U__d1, U__d0, P[40]);
  U4DPPG_25_8 U25 (P[42], O_R[41], IN1_R[25], U__d1, U__d0, P[41]);
  U4DPPG_26_8 U26 (P[43], O_R[42], IN1_R[26], U__d1, U__d0, P[42]);
  U4DPPG_27_8 U27 (P[44], O_R[43], IN1_R[27], U__d1, U__d0, P[43]);
  U4DPPG_28_8 U28 (P[45], O_R[44], IN1_R[28], U__d1, U__d0, P[44]);
  U4DPPG_29_8 U29 (P[46], O_R[45], IN1_R[29], U__d1, U__d0, P[45]);
  U4DPPG_30_8 U30 (P[47], O_R[46], IN1_R[30], U__d1, U__d0, P[46]);
  U4DPPG_31_8 U31 (P[48], O_R[47], IN1_R[31], U__d1, U__d0, P[47]);
  U4DPPG_32_8 U32 (P[49], O_R[48], IN1_R[32], U__d1, U__d0, P[48]);
  U4DPPG_33_8 U33 (P[50], O_R[49], IN1_R[33], U__d1, U__d0, P[49]);
  U4DPPG_34_8 U34 (P[51], O_R[50], IN1_R[34], U__d1, U__d0, P[50]);
  U4DPPG_35_8 U35 (P[52], O_R[51], IN1_R[35], U__d1, U__d0, P[51]);
  U4DPPG_36_8 U36 (P[53], O_R[52], IN1_R[36], U__d1, U__d0, P[52]);
  U4DPPG_37_8 U37 (P[54], O_R[53], IN1_R[37], U__d1, U__d0, P[53]);
  U4DPPG_38_8 U38 (P[55], O_R[54], IN1_R[38], U__d1, U__d0, P[54]);
  U4DPPG_39_8 U39 (P[56], O_R[55], IN1_R[39], U__d1, U__d0, P[55]);
  U4DPPG_40_8 U40 (P[57], O_R[56], IN1_R[40], U__d1, U__d0, P[56]);
  U4DPPG_41_8 U41 (P[58], O_R[57], IN1_R[41], U__d1, U__d0, P[57]);
  U4DPPG_42_8 U42 (P[59], O_R[58], IN1_R[42], U__d1, U__d0, P[58]);
  U4DPPG_43_8 U43 (P[60], O_R[59], IN1_R[43], U__d1, U__d0, P[59]);
  U4DPPG_44_8 U44 (P[61], O_R[60], IN1_R[44], U__d1, U__d0, P[60]);
  U4DPPG_45_8 U45 (P[62], O_R[61], IN1_R[45], U__d1, U__d0, P[61]);
  U4DPPG_46_8 U46 (P[63], O_R[62], IN1_R[46], U__d1, U__d0, P[62]);
  U4DPPG_47_8 U47 (P[64], O_R[63], IN1_R[47], U__d1, U__d0, P[63]);
  U4DPPG_48_8 U48 (P[65], O_R[64], IN1_R[48], U__d1, U__d0, P[64]);
  U4DPPG_49_8 U49 (P[66], O_R[65], IN1_R[49], U__d1, U__d0, P[65]);
  U4DPPG_50_8 U50 (P[67], O_R[66], IN1_R[50], U__d1, U__d0, P[66]);
  U4DPPG_51_8 U51 (P[68], O_R[67], IN1_R[51], U__d1, U__d0, P[67]);
  U4DPPG_52_8 U52 (P[69], O_R[68], IN1_R[52], U__d1, U__d0, P[68]);
  U4DPPG_53_8 U53 (P[70], O_R[69], IN1_R[53], U__d1, U__d0, P[69]);
  U4DPPG_54_8 U54 (P[71], O_R[70], IN1_R[54], U__d1, U__d0, P[70]);
  U4DPPG_55_8 U55 (P[72], O_R[71], IN1_R[55], U__d1, U__d0, P[71]);
  U4DPPG_56_8 U56 (P[73], O_R[72], IN1_R[56], U__d1, U__d0, P[72]);
  U4DPPG_57_8 U57 (P[74], O_R[73], IN1_R[57], U__d1, U__d0, P[73]);
  U4DPPG_58_8 U58 (P[75], O_R[74], IN1_R[58], U__d1, U__d0, P[74]);
  U4DPPG_59_8 U59 (P[76], O_R[75], IN1_R[59], U__d1, U__d0, P[75]);
  U4DPPG_60_8 U60 (P[77], O_R[76], IN1_R[60], U__d1, U__d0, P[76]);
  U4DPPG_61_8 U61 (P[78], O_R[77], IN1_R[61], U__d1, U__d0, P[77]);
  U4DPPG_62_8 U62 (P[79], O_R[78], IN1_R[62], U__d1, U__d0, P[78]);
  U4DPPGH_63_8 U63 (O_T, O_R[79], IN1_T, U__d1, U__d0, P[79]);
endmodule

module TCU4VPPG_63_0_9 (O_T, O_R, IN1_T, IN1_R, U__d1, U__d0);
  output [81:18] O_R;
  output O_T;
  input [62:0] IN1_R;
  input IN1_T;
  input U__d1, U__d0;
  wire [81:19] P;
  U4DPPGL_0_9 U0 (P[19], O_R[18], IN1_R[0], U__d1, U__d0);
  U4DPPG_1_9 U1 (P[20], O_R[19], IN1_R[1], U__d1, U__d0, P[19]);
  U4DPPG_2_9 U2 (P[21], O_R[20], IN1_R[2], U__d1, U__d0, P[20]);
  U4DPPG_3_9 U3 (P[22], O_R[21], IN1_R[3], U__d1, U__d0, P[21]);
  U4DPPG_4_9 U4 (P[23], O_R[22], IN1_R[4], U__d1, U__d0, P[22]);
  U4DPPG_5_9 U5 (P[24], O_R[23], IN1_R[5], U__d1, U__d0, P[23]);
  U4DPPG_6_9 U6 (P[25], O_R[24], IN1_R[6], U__d1, U__d0, P[24]);
  U4DPPG_7_9 U7 (P[26], O_R[25], IN1_R[7], U__d1, U__d0, P[25]);
  U4DPPG_8_9 U8 (P[27], O_R[26], IN1_R[8], U__d1, U__d0, P[26]);
  U4DPPG_9_9 U9 (P[28], O_R[27], IN1_R[9], U__d1, U__d0, P[27]);
  U4DPPG_10_9 U10 (P[29], O_R[28], IN1_R[10], U__d1, U__d0, P[28]);
  U4DPPG_11_9 U11 (P[30], O_R[29], IN1_R[11], U__d1, U__d0, P[29]);
  U4DPPG_12_9 U12 (P[31], O_R[30], IN1_R[12], U__d1, U__d0, P[30]);
  U4DPPG_13_9 U13 (P[32], O_R[31], IN1_R[13], U__d1, U__d0, P[31]);
  U4DPPG_14_9 U14 (P[33], O_R[32], IN1_R[14], U__d1, U__d0, P[32]);
  U4DPPG_15_9 U15 (P[34], O_R[33], IN1_R[15], U__d1, U__d0, P[33]);
  U4DPPG_16_9 U16 (P[35], O_R[34], IN1_R[16], U__d1, U__d0, P[34]);
  U4DPPG_17_9 U17 (P[36], O_R[35], IN1_R[17], U__d1, U__d0, P[35]);
  U4DPPG_18_9 U18 (P[37], O_R[36], IN1_R[18], U__d1, U__d0, P[36]);
  U4DPPG_19_9 U19 (P[38], O_R[37], IN1_R[19], U__d1, U__d0, P[37]);
  U4DPPG_20_9 U20 (P[39], O_R[38], IN1_R[20], U__d1, U__d0, P[38]);
  U4DPPG_21_9 U21 (P[40], O_R[39], IN1_R[21], U__d1, U__d0, P[39]);
  U4DPPG_22_9 U22 (P[41], O_R[40], IN1_R[22], U__d1, U__d0, P[40]);
  U4DPPG_23_9 U23 (P[42], O_R[41], IN1_R[23], U__d1, U__d0, P[41]);
  U4DPPG_24_9 U24 (P[43], O_R[42], IN1_R[24], U__d1, U__d0, P[42]);
  U4DPPG_25_9 U25 (P[44], O_R[43], IN1_R[25], U__d1, U__d0, P[43]);
  U4DPPG_26_9 U26 (P[45], O_R[44], IN1_R[26], U__d1, U__d0, P[44]);
  U4DPPG_27_9 U27 (P[46], O_R[45], IN1_R[27], U__d1, U__d0, P[45]);
  U4DPPG_28_9 U28 (P[47], O_R[46], IN1_R[28], U__d1, U__d0, P[46]);
  U4DPPG_29_9 U29 (P[48], O_R[47], IN1_R[29], U__d1, U__d0, P[47]);
  U4DPPG_30_9 U30 (P[49], O_R[48], IN1_R[30], U__d1, U__d0, P[48]);
  U4DPPG_31_9 U31 (P[50], O_R[49], IN1_R[31], U__d1, U__d0, P[49]);
  U4DPPG_32_9 U32 (P[51], O_R[50], IN1_R[32], U__d1, U__d0, P[50]);
  U4DPPG_33_9 U33 (P[52], O_R[51], IN1_R[33], U__d1, U__d0, P[51]);
  U4DPPG_34_9 U34 (P[53], O_R[52], IN1_R[34], U__d1, U__d0, P[52]);
  U4DPPG_35_9 U35 (P[54], O_R[53], IN1_R[35], U__d1, U__d0, P[53]);
  U4DPPG_36_9 U36 (P[55], O_R[54], IN1_R[36], U__d1, U__d0, P[54]);
  U4DPPG_37_9 U37 (P[56], O_R[55], IN1_R[37], U__d1, U__d0, P[55]);
  U4DPPG_38_9 U38 (P[57], O_R[56], IN1_R[38], U__d1, U__d0, P[56]);
  U4DPPG_39_9 U39 (P[58], O_R[57], IN1_R[39], U__d1, U__d0, P[57]);
  U4DPPG_40_9 U40 (P[59], O_R[58], IN1_R[40], U__d1, U__d0, P[58]);
  U4DPPG_41_9 U41 (P[60], O_R[59], IN1_R[41], U__d1, U__d0, P[59]);
  U4DPPG_42_9 U42 (P[61], O_R[60], IN1_R[42], U__d1, U__d0, P[60]);
  U4DPPG_43_9 U43 (P[62], O_R[61], IN1_R[43], U__d1, U__d0, P[61]);
  U4DPPG_44_9 U44 (P[63], O_R[62], IN1_R[44], U__d1, U__d0, P[62]);
  U4DPPG_45_9 U45 (P[64], O_R[63], IN1_R[45], U__d1, U__d0, P[63]);
  U4DPPG_46_9 U46 (P[65], O_R[64], IN1_R[46], U__d1, U__d0, P[64]);
  U4DPPG_47_9 U47 (P[66], O_R[65], IN1_R[47], U__d1, U__d0, P[65]);
  U4DPPG_48_9 U48 (P[67], O_R[66], IN1_R[48], U__d1, U__d0, P[66]);
  U4DPPG_49_9 U49 (P[68], O_R[67], IN1_R[49], U__d1, U__d0, P[67]);
  U4DPPG_50_9 U50 (P[69], O_R[68], IN1_R[50], U__d1, U__d0, P[68]);
  U4DPPG_51_9 U51 (P[70], O_R[69], IN1_R[51], U__d1, U__d0, P[69]);
  U4DPPG_52_9 U52 (P[71], O_R[70], IN1_R[52], U__d1, U__d0, P[70]);
  U4DPPG_53_9 U53 (P[72], O_R[71], IN1_R[53], U__d1, U__d0, P[71]);
  U4DPPG_54_9 U54 (P[73], O_R[72], IN1_R[54], U__d1, U__d0, P[72]);
  U4DPPG_55_9 U55 (P[74], O_R[73], IN1_R[55], U__d1, U__d0, P[73]);
  U4DPPG_56_9 U56 (P[75], O_R[74], IN1_R[56], U__d1, U__d0, P[74]);
  U4DPPG_57_9 U57 (P[76], O_R[75], IN1_R[57], U__d1, U__d0, P[75]);
  U4DPPG_58_9 U58 (P[77], O_R[76], IN1_R[58], U__d1, U__d0, P[76]);
  U4DPPG_59_9 U59 (P[78], O_R[77], IN1_R[59], U__d1, U__d0, P[77]);
  U4DPPG_60_9 U60 (P[79], O_R[78], IN1_R[60], U__d1, U__d0, P[78]);
  U4DPPG_61_9 U61 (P[80], O_R[79], IN1_R[61], U__d1, U__d0, P[79]);
  U4DPPG_62_9 U62 (P[81], O_R[80], IN1_R[62], U__d1, U__d0, P[80]);
  U4DPPGH_63_9 U63 (O_T, O_R[81], IN1_T, U__d1, U__d0, P[81]);
endmodule

module TUBWCON_100_36 (O, I_T, I_R, S);
  output [100:36] O;
  input [99:36] I_R;
  input I_T;
  input S;
  BWCPP_36 U0 (O[36], I_R[36], S);
  BWCPP_37 U1 (O[37], I_R[37], S);
  BWCPP_38 U2 (O[38], I_R[38], S);
  BWCPP_39 U3 (O[39], I_R[39], S);
  BWCPP_40 U4 (O[40], I_R[40], S);
  BWCPP_41 U5 (O[41], I_R[41], S);
  BWCPP_42 U6 (O[42], I_R[42], S);
  BWCPP_43 U7 (O[43], I_R[43], S);
  BWCPP_44 U8 (O[44], I_R[44], S);
  BWCPP_45 U9 (O[45], I_R[45], S);
  BWCPP_46 U10 (O[46], I_R[46], S);
  BWCPP_47 U11 (O[47], I_R[47], S);
  BWCPP_48 U12 (O[48], I_R[48], S);
  BWCPP_49 U13 (O[49], I_R[49], S);
  BWCPP_50 U14 (O[50], I_R[50], S);
  BWCPP_51 U15 (O[51], I_R[51], S);
  BWCPP_52 U16 (O[52], I_R[52], S);
  BWCPP_53 U17 (O[53], I_R[53], S);
  BWCPP_54 U18 (O[54], I_R[54], S);
  BWCPP_55 U19 (O[55], I_R[55], S);
  BWCPP_56 U20 (O[56], I_R[56], S);
  BWCPP_57 U21 (O[57], I_R[57], S);
  BWCPP_58 U22 (O[58], I_R[58], S);
  BWCPP_59 U23 (O[59], I_R[59], S);
  BWCPP_60 U24 (O[60], I_R[60], S);
  BWCPP_61 U25 (O[61], I_R[61], S);
  BWCPP_62 U26 (O[62], I_R[62], S);
  BWCPP_63 U27 (O[63], I_R[63], S);
  BWCPP_64 U28 (O[64], I_R[64], S);
  BWCPP_65 U29 (O[65], I_R[65], S);
  BWCPP_66 U30 (O[66], I_R[66], S);
  BWCPP_67 U31 (O[67], I_R[67], S);
  BWCPP_68 U32 (O[68], I_R[68], S);
  BWCPP_69 U33 (O[69], I_R[69], S);
  BWCPP_70 U34 (O[70], I_R[70], S);
  BWCPP_71 U35 (O[71], I_R[71], S);
  BWCPP_72 U36 (O[72], I_R[72], S);
  BWCPP_73 U37 (O[73], I_R[73], S);
  BWCPP_74 U38 (O[74], I_R[74], S);
  BWCPP_75 U39 (O[75], I_R[75], S);
  BWCPP_76 U40 (O[76], I_R[76], S);
  BWCPP_77 U41 (O[77], I_R[77], S);
  BWCPP_78 U42 (O[78], I_R[78], S);
  BWCPP_79 U43 (O[79], I_R[79], S);
  BWCPP_80 U44 (O[80], I_R[80], S);
  BWCPP_81 U45 (O[81], I_R[81], S);
  BWCPP_82 U46 (O[82], I_R[82], S);
  BWCPP_83 U47 (O[83], I_R[83], S);
  BWCPP_84 U48 (O[84], I_R[84], S);
  BWCPP_85 U49 (O[85], I_R[85], S);
  BWCPP_86 U50 (O[86], I_R[86], S);
  BWCPP_87 U51 (O[87], I_R[87], S);
  BWCPP_88 U52 (O[88], I_R[88], S);
  BWCPP_89 U53 (O[89], I_R[89], S);
  BWCPP_90 U54 (O[90], I_R[90], S);
  BWCPP_91 U55 (O[91], I_R[91], S);
  BWCPP_92 U56 (O[92], I_R[92], S);
  BWCPP_93 U57 (O[93], I_R[93], S);
  BWCPP_94 U58 (O[94], I_R[94], S);
  BWCPP_95 U59 (O[95], I_R[95], S);
  BWCPP_96 U60 (O[96], I_R[96], S);
  BWCPP_97 U61 (O[97], I_R[97], S);
  BWCPP_98 U62 (O[98], I_R[98], S);
  BWCPP_99 U63 (O[99], I_R[99], S);
  BWCNP_100 U64 (O[100], I_T, S);
endmodule

module TUBWCON_102_38 (O, I_T, I_R, S);
  output [102:38] O;
  input [101:38] I_R;
  input I_T;
  input S;
  BWCPP_38 U0 (O[38], I_R[38], S);
  BWCPP_39 U1 (O[39], I_R[39], S);
  BWCPP_40 U2 (O[40], I_R[40], S);
  BWCPP_41 U3 (O[41], I_R[41], S);
  BWCPP_42 U4 (O[42], I_R[42], S);
  BWCPP_43 U5 (O[43], I_R[43], S);
  BWCPP_44 U6 (O[44], I_R[44], S);
  BWCPP_45 U7 (O[45], I_R[45], S);
  BWCPP_46 U8 (O[46], I_R[46], S);
  BWCPP_47 U9 (O[47], I_R[47], S);
  BWCPP_48 U10 (O[48], I_R[48], S);
  BWCPP_49 U11 (O[49], I_R[49], S);
  BWCPP_50 U12 (O[50], I_R[50], S);
  BWCPP_51 U13 (O[51], I_R[51], S);
  BWCPP_52 U14 (O[52], I_R[52], S);
  BWCPP_53 U15 (O[53], I_R[53], S);
  BWCPP_54 U16 (O[54], I_R[54], S);
  BWCPP_55 U17 (O[55], I_R[55], S);
  BWCPP_56 U18 (O[56], I_R[56], S);
  BWCPP_57 U19 (O[57], I_R[57], S);
  BWCPP_58 U20 (O[58], I_R[58], S);
  BWCPP_59 U21 (O[59], I_R[59], S);
  BWCPP_60 U22 (O[60], I_R[60], S);
  BWCPP_61 U23 (O[61], I_R[61], S);
  BWCPP_62 U24 (O[62], I_R[62], S);
  BWCPP_63 U25 (O[63], I_R[63], S);
  BWCPP_64 U26 (O[64], I_R[64], S);
  BWCPP_65 U27 (O[65], I_R[65], S);
  BWCPP_66 U28 (O[66], I_R[66], S);
  BWCPP_67 U29 (O[67], I_R[67], S);
  BWCPP_68 U30 (O[68], I_R[68], S);
  BWCPP_69 U31 (O[69], I_R[69], S);
  BWCPP_70 U32 (O[70], I_R[70], S);
  BWCPP_71 U33 (O[71], I_R[71], S);
  BWCPP_72 U34 (O[72], I_R[72], S);
  BWCPP_73 U35 (O[73], I_R[73], S);
  BWCPP_74 U36 (O[74], I_R[74], S);
  BWCPP_75 U37 (O[75], I_R[75], S);
  BWCPP_76 U38 (O[76], I_R[76], S);
  BWCPP_77 U39 (O[77], I_R[77], S);
  BWCPP_78 U40 (O[78], I_R[78], S);
  BWCPP_79 U41 (O[79], I_R[79], S);
  BWCPP_80 U42 (O[80], I_R[80], S);
  BWCPP_81 U43 (O[81], I_R[81], S);
  BWCPP_82 U44 (O[82], I_R[82], S);
  BWCPP_83 U45 (O[83], I_R[83], S);
  BWCPP_84 U46 (O[84], I_R[84], S);
  BWCPP_85 U47 (O[85], I_R[85], S);
  BWCPP_86 U48 (O[86], I_R[86], S);
  BWCPP_87 U49 (O[87], I_R[87], S);
  BWCPP_88 U50 (O[88], I_R[88], S);
  BWCPP_89 U51 (O[89], I_R[89], S);
  BWCPP_90 U52 (O[90], I_R[90], S);
  BWCPP_91 U53 (O[91], I_R[91], S);
  BWCPP_92 U54 (O[92], I_R[92], S);
  BWCPP_93 U55 (O[93], I_R[93], S);
  BWCPP_94 U56 (O[94], I_R[94], S);
  BWCPP_95 U57 (O[95], I_R[95], S);
  BWCPP_96 U58 (O[96], I_R[96], S);
  BWCPP_97 U59 (O[97], I_R[97], S);
  BWCPP_98 U60 (O[98], I_R[98], S);
  BWCPP_99 U61 (O[99], I_R[99], S);
  BWCPP_100 U62 (O[100], I_R[100], S);
  BWCPP_101 U63 (O[101], I_R[101], S);
  BWCNP_102 U64 (O[102], I_T, S);
endmodule

module TUBWCON_104_40 (O, I_T, I_R, S);
  output [104:40] O;
  input [103:40] I_R;
  input I_T;
  input S;
  BWCPP_40 U0 (O[40], I_R[40], S);
  BWCPP_41 U1 (O[41], I_R[41], S);
  BWCPP_42 U2 (O[42], I_R[42], S);
  BWCPP_43 U3 (O[43], I_R[43], S);
  BWCPP_44 U4 (O[44], I_R[44], S);
  BWCPP_45 U5 (O[45], I_R[45], S);
  BWCPP_46 U6 (O[46], I_R[46], S);
  BWCPP_47 U7 (O[47], I_R[47], S);
  BWCPP_48 U8 (O[48], I_R[48], S);
  BWCPP_49 U9 (O[49], I_R[49], S);
  BWCPP_50 U10 (O[50], I_R[50], S);
  BWCPP_51 U11 (O[51], I_R[51], S);
  BWCPP_52 U12 (O[52], I_R[52], S);
  BWCPP_53 U13 (O[53], I_R[53], S);
  BWCPP_54 U14 (O[54], I_R[54], S);
  BWCPP_55 U15 (O[55], I_R[55], S);
  BWCPP_56 U16 (O[56], I_R[56], S);
  BWCPP_57 U17 (O[57], I_R[57], S);
  BWCPP_58 U18 (O[58], I_R[58], S);
  BWCPP_59 U19 (O[59], I_R[59], S);
  BWCPP_60 U20 (O[60], I_R[60], S);
  BWCPP_61 U21 (O[61], I_R[61], S);
  BWCPP_62 U22 (O[62], I_R[62], S);
  BWCPP_63 U23 (O[63], I_R[63], S);
  BWCPP_64 U24 (O[64], I_R[64], S);
  BWCPP_65 U25 (O[65], I_R[65], S);
  BWCPP_66 U26 (O[66], I_R[66], S);
  BWCPP_67 U27 (O[67], I_R[67], S);
  BWCPP_68 U28 (O[68], I_R[68], S);
  BWCPP_69 U29 (O[69], I_R[69], S);
  BWCPP_70 U30 (O[70], I_R[70], S);
  BWCPP_71 U31 (O[71], I_R[71], S);
  BWCPP_72 U32 (O[72], I_R[72], S);
  BWCPP_73 U33 (O[73], I_R[73], S);
  BWCPP_74 U34 (O[74], I_R[74], S);
  BWCPP_75 U35 (O[75], I_R[75], S);
  BWCPP_76 U36 (O[76], I_R[76], S);
  BWCPP_77 U37 (O[77], I_R[77], S);
  BWCPP_78 U38 (O[78], I_R[78], S);
  BWCPP_79 U39 (O[79], I_R[79], S);
  BWCPP_80 U40 (O[80], I_R[80], S);
  BWCPP_81 U41 (O[81], I_R[81], S);
  BWCPP_82 U42 (O[82], I_R[82], S);
  BWCPP_83 U43 (O[83], I_R[83], S);
  BWCPP_84 U44 (O[84], I_R[84], S);
  BWCPP_85 U45 (O[85], I_R[85], S);
  BWCPP_86 U46 (O[86], I_R[86], S);
  BWCPP_87 U47 (O[87], I_R[87], S);
  BWCPP_88 U48 (O[88], I_R[88], S);
  BWCPP_89 U49 (O[89], I_R[89], S);
  BWCPP_90 U50 (O[90], I_R[90], S);
  BWCPP_91 U51 (O[91], I_R[91], S);
  BWCPP_92 U52 (O[92], I_R[92], S);
  BWCPP_93 U53 (O[93], I_R[93], S);
  BWCPP_94 U54 (O[94], I_R[94], S);
  BWCPP_95 U55 (O[95], I_R[95], S);
  BWCPP_96 U56 (O[96], I_R[96], S);
  BWCPP_97 U57 (O[97], I_R[97], S);
  BWCPP_98 U58 (O[98], I_R[98], S);
  BWCPP_99 U59 (O[99], I_R[99], S);
  BWCPP_100 U60 (O[100], I_R[100], S);
  BWCPP_101 U61 (O[101], I_R[101], S);
  BWCPP_102 U62 (O[102], I_R[102], S);
  BWCPP_103 U63 (O[103], I_R[103], S);
  BWCNP_104 U64 (O[104], I_T, S);
endmodule

module TUBWCON_106_42 (O, I_T, I_R, S);
  output [106:42] O;
  input [105:42] I_R;
  input I_T;
  input S;
  BWCPP_42 U0 (O[42], I_R[42], S);
  BWCPP_43 U1 (O[43], I_R[43], S);
  BWCPP_44 U2 (O[44], I_R[44], S);
  BWCPP_45 U3 (O[45], I_R[45], S);
  BWCPP_46 U4 (O[46], I_R[46], S);
  BWCPP_47 U5 (O[47], I_R[47], S);
  BWCPP_48 U6 (O[48], I_R[48], S);
  BWCPP_49 U7 (O[49], I_R[49], S);
  BWCPP_50 U8 (O[50], I_R[50], S);
  BWCPP_51 U9 (O[51], I_R[51], S);
  BWCPP_52 U10 (O[52], I_R[52], S);
  BWCPP_53 U11 (O[53], I_R[53], S);
  BWCPP_54 U12 (O[54], I_R[54], S);
  BWCPP_55 U13 (O[55], I_R[55], S);
  BWCPP_56 U14 (O[56], I_R[56], S);
  BWCPP_57 U15 (O[57], I_R[57], S);
  BWCPP_58 U16 (O[58], I_R[58], S);
  BWCPP_59 U17 (O[59], I_R[59], S);
  BWCPP_60 U18 (O[60], I_R[60], S);
  BWCPP_61 U19 (O[61], I_R[61], S);
  BWCPP_62 U20 (O[62], I_R[62], S);
  BWCPP_63 U21 (O[63], I_R[63], S);
  BWCPP_64 U22 (O[64], I_R[64], S);
  BWCPP_65 U23 (O[65], I_R[65], S);
  BWCPP_66 U24 (O[66], I_R[66], S);
  BWCPP_67 U25 (O[67], I_R[67], S);
  BWCPP_68 U26 (O[68], I_R[68], S);
  BWCPP_69 U27 (O[69], I_R[69], S);
  BWCPP_70 U28 (O[70], I_R[70], S);
  BWCPP_71 U29 (O[71], I_R[71], S);
  BWCPP_72 U30 (O[72], I_R[72], S);
  BWCPP_73 U31 (O[73], I_R[73], S);
  BWCPP_74 U32 (O[74], I_R[74], S);
  BWCPP_75 U33 (O[75], I_R[75], S);
  BWCPP_76 U34 (O[76], I_R[76], S);
  BWCPP_77 U35 (O[77], I_R[77], S);
  BWCPP_78 U36 (O[78], I_R[78], S);
  BWCPP_79 U37 (O[79], I_R[79], S);
  BWCPP_80 U38 (O[80], I_R[80], S);
  BWCPP_81 U39 (O[81], I_R[81], S);
  BWCPP_82 U40 (O[82], I_R[82], S);
  BWCPP_83 U41 (O[83], I_R[83], S);
  BWCPP_84 U42 (O[84], I_R[84], S);
  BWCPP_85 U43 (O[85], I_R[85], S);
  BWCPP_86 U44 (O[86], I_R[86], S);
  BWCPP_87 U45 (O[87], I_R[87], S);
  BWCPP_88 U46 (O[88], I_R[88], S);
  BWCPP_89 U47 (O[89], I_R[89], S);
  BWCPP_90 U48 (O[90], I_R[90], S);
  BWCPP_91 U49 (O[91], I_R[91], S);
  BWCPP_92 U50 (O[92], I_R[92], S);
  BWCPP_93 U51 (O[93], I_R[93], S);
  BWCPP_94 U52 (O[94], I_R[94], S);
  BWCPP_95 U53 (O[95], I_R[95], S);
  BWCPP_96 U54 (O[96], I_R[96], S);
  BWCPP_97 U55 (O[97], I_R[97], S);
  BWCPP_98 U56 (O[98], I_R[98], S);
  BWCPP_99 U57 (O[99], I_R[99], S);
  BWCPP_100 U58 (O[100], I_R[100], S);
  BWCPP_101 U59 (O[101], I_R[101], S);
  BWCPP_102 U60 (O[102], I_R[102], S);
  BWCPP_103 U61 (O[103], I_R[103], S);
  BWCPP_104 U62 (O[104], I_R[104], S);
  BWCPP_105 U63 (O[105], I_R[105], S);
  BWCNP_106 U64 (O[106], I_T, S);
endmodule

module TUBWCON_108_44 (O, I_T, I_R, S);
  output [108:44] O;
  input [107:44] I_R;
  input I_T;
  input S;
  BWCPP_44 U0 (O[44], I_R[44], S);
  BWCPP_45 U1 (O[45], I_R[45], S);
  BWCPP_46 U2 (O[46], I_R[46], S);
  BWCPP_47 U3 (O[47], I_R[47], S);
  BWCPP_48 U4 (O[48], I_R[48], S);
  BWCPP_49 U5 (O[49], I_R[49], S);
  BWCPP_50 U6 (O[50], I_R[50], S);
  BWCPP_51 U7 (O[51], I_R[51], S);
  BWCPP_52 U8 (O[52], I_R[52], S);
  BWCPP_53 U9 (O[53], I_R[53], S);
  BWCPP_54 U10 (O[54], I_R[54], S);
  BWCPP_55 U11 (O[55], I_R[55], S);
  BWCPP_56 U12 (O[56], I_R[56], S);
  BWCPP_57 U13 (O[57], I_R[57], S);
  BWCPP_58 U14 (O[58], I_R[58], S);
  BWCPP_59 U15 (O[59], I_R[59], S);
  BWCPP_60 U16 (O[60], I_R[60], S);
  BWCPP_61 U17 (O[61], I_R[61], S);
  BWCPP_62 U18 (O[62], I_R[62], S);
  BWCPP_63 U19 (O[63], I_R[63], S);
  BWCPP_64 U20 (O[64], I_R[64], S);
  BWCPP_65 U21 (O[65], I_R[65], S);
  BWCPP_66 U22 (O[66], I_R[66], S);
  BWCPP_67 U23 (O[67], I_R[67], S);
  BWCPP_68 U24 (O[68], I_R[68], S);
  BWCPP_69 U25 (O[69], I_R[69], S);
  BWCPP_70 U26 (O[70], I_R[70], S);
  BWCPP_71 U27 (O[71], I_R[71], S);
  BWCPP_72 U28 (O[72], I_R[72], S);
  BWCPP_73 U29 (O[73], I_R[73], S);
  BWCPP_74 U30 (O[74], I_R[74], S);
  BWCPP_75 U31 (O[75], I_R[75], S);
  BWCPP_76 U32 (O[76], I_R[76], S);
  BWCPP_77 U33 (O[77], I_R[77], S);
  BWCPP_78 U34 (O[78], I_R[78], S);
  BWCPP_79 U35 (O[79], I_R[79], S);
  BWCPP_80 U36 (O[80], I_R[80], S);
  BWCPP_81 U37 (O[81], I_R[81], S);
  BWCPP_82 U38 (O[82], I_R[82], S);
  BWCPP_83 U39 (O[83], I_R[83], S);
  BWCPP_84 U40 (O[84], I_R[84], S);
  BWCPP_85 U41 (O[85], I_R[85], S);
  BWCPP_86 U42 (O[86], I_R[86], S);
  BWCPP_87 U43 (O[87], I_R[87], S);
  BWCPP_88 U44 (O[88], I_R[88], S);
  BWCPP_89 U45 (O[89], I_R[89], S);
  BWCPP_90 U46 (O[90], I_R[90], S);
  BWCPP_91 U47 (O[91], I_R[91], S);
  BWCPP_92 U48 (O[92], I_R[92], S);
  BWCPP_93 U49 (O[93], I_R[93], S);
  BWCPP_94 U50 (O[94], I_R[94], S);
  BWCPP_95 U51 (O[95], I_R[95], S);
  BWCPP_96 U52 (O[96], I_R[96], S);
  BWCPP_97 U53 (O[97], I_R[97], S);
  BWCPP_98 U54 (O[98], I_R[98], S);
  BWCPP_99 U55 (O[99], I_R[99], S);
  BWCPP_100 U56 (O[100], I_R[100], S);
  BWCPP_101 U57 (O[101], I_R[101], S);
  BWCPP_102 U58 (O[102], I_R[102], S);
  BWCPP_103 U59 (O[103], I_R[103], S);
  BWCPP_104 U60 (O[104], I_R[104], S);
  BWCPP_105 U61 (O[105], I_R[105], S);
  BWCPP_106 U62 (O[106], I_R[106], S);
  BWCPP_107 U63 (O[107], I_R[107], S);
  BWCNP_108 U64 (O[108], I_T, S);
endmodule

module TUBWCON_110_46 (O, I_T, I_R, S);
  output [110:46] O;
  input [109:46] I_R;
  input I_T;
  input S;
  BWCPP_46 U0 (O[46], I_R[46], S);
  BWCPP_47 U1 (O[47], I_R[47], S);
  BWCPP_48 U2 (O[48], I_R[48], S);
  BWCPP_49 U3 (O[49], I_R[49], S);
  BWCPP_50 U4 (O[50], I_R[50], S);
  BWCPP_51 U5 (O[51], I_R[51], S);
  BWCPP_52 U6 (O[52], I_R[52], S);
  BWCPP_53 U7 (O[53], I_R[53], S);
  BWCPP_54 U8 (O[54], I_R[54], S);
  BWCPP_55 U9 (O[55], I_R[55], S);
  BWCPP_56 U10 (O[56], I_R[56], S);
  BWCPP_57 U11 (O[57], I_R[57], S);
  BWCPP_58 U12 (O[58], I_R[58], S);
  BWCPP_59 U13 (O[59], I_R[59], S);
  BWCPP_60 U14 (O[60], I_R[60], S);
  BWCPP_61 U15 (O[61], I_R[61], S);
  BWCPP_62 U16 (O[62], I_R[62], S);
  BWCPP_63 U17 (O[63], I_R[63], S);
  BWCPP_64 U18 (O[64], I_R[64], S);
  BWCPP_65 U19 (O[65], I_R[65], S);
  BWCPP_66 U20 (O[66], I_R[66], S);
  BWCPP_67 U21 (O[67], I_R[67], S);
  BWCPP_68 U22 (O[68], I_R[68], S);
  BWCPP_69 U23 (O[69], I_R[69], S);
  BWCPP_70 U24 (O[70], I_R[70], S);
  BWCPP_71 U25 (O[71], I_R[71], S);
  BWCPP_72 U26 (O[72], I_R[72], S);
  BWCPP_73 U27 (O[73], I_R[73], S);
  BWCPP_74 U28 (O[74], I_R[74], S);
  BWCPP_75 U29 (O[75], I_R[75], S);
  BWCPP_76 U30 (O[76], I_R[76], S);
  BWCPP_77 U31 (O[77], I_R[77], S);
  BWCPP_78 U32 (O[78], I_R[78], S);
  BWCPP_79 U33 (O[79], I_R[79], S);
  BWCPP_80 U34 (O[80], I_R[80], S);
  BWCPP_81 U35 (O[81], I_R[81], S);
  BWCPP_82 U36 (O[82], I_R[82], S);
  BWCPP_83 U37 (O[83], I_R[83], S);
  BWCPP_84 U38 (O[84], I_R[84], S);
  BWCPP_85 U39 (O[85], I_R[85], S);
  BWCPP_86 U40 (O[86], I_R[86], S);
  BWCPP_87 U41 (O[87], I_R[87], S);
  BWCPP_88 U42 (O[88], I_R[88], S);
  BWCPP_89 U43 (O[89], I_R[89], S);
  BWCPP_90 U44 (O[90], I_R[90], S);
  BWCPP_91 U45 (O[91], I_R[91], S);
  BWCPP_92 U46 (O[92], I_R[92], S);
  BWCPP_93 U47 (O[93], I_R[93], S);
  BWCPP_94 U48 (O[94], I_R[94], S);
  BWCPP_95 U49 (O[95], I_R[95], S);
  BWCPP_96 U50 (O[96], I_R[96], S);
  BWCPP_97 U51 (O[97], I_R[97], S);
  BWCPP_98 U52 (O[98], I_R[98], S);
  BWCPP_99 U53 (O[99], I_R[99], S);
  BWCPP_100 U54 (O[100], I_R[100], S);
  BWCPP_101 U55 (O[101], I_R[101], S);
  BWCPP_102 U56 (O[102], I_R[102], S);
  BWCPP_103 U57 (O[103], I_R[103], S);
  BWCPP_104 U58 (O[104], I_R[104], S);
  BWCPP_105 U59 (O[105], I_R[105], S);
  BWCPP_106 U60 (O[106], I_R[106], S);
  BWCPP_107 U61 (O[107], I_R[107], S);
  BWCPP_108 U62 (O[108], I_R[108], S);
  BWCPP_109 U63 (O[109], I_R[109], S);
  BWCNP_110 U64 (O[110], I_T, S);
endmodule

module TUBWCON_112_48 (O, I_T, I_R, S);
  output [112:48] O;
  input [111:48] I_R;
  input I_T;
  input S;
  BWCPP_48 U0 (O[48], I_R[48], S);
  BWCPP_49 U1 (O[49], I_R[49], S);
  BWCPP_50 U2 (O[50], I_R[50], S);
  BWCPP_51 U3 (O[51], I_R[51], S);
  BWCPP_52 U4 (O[52], I_R[52], S);
  BWCPP_53 U5 (O[53], I_R[53], S);
  BWCPP_54 U6 (O[54], I_R[54], S);
  BWCPP_55 U7 (O[55], I_R[55], S);
  BWCPP_56 U8 (O[56], I_R[56], S);
  BWCPP_57 U9 (O[57], I_R[57], S);
  BWCPP_58 U10 (O[58], I_R[58], S);
  BWCPP_59 U11 (O[59], I_R[59], S);
  BWCPP_60 U12 (O[60], I_R[60], S);
  BWCPP_61 U13 (O[61], I_R[61], S);
  BWCPP_62 U14 (O[62], I_R[62], S);
  BWCPP_63 U15 (O[63], I_R[63], S);
  BWCPP_64 U16 (O[64], I_R[64], S);
  BWCPP_65 U17 (O[65], I_R[65], S);
  BWCPP_66 U18 (O[66], I_R[66], S);
  BWCPP_67 U19 (O[67], I_R[67], S);
  BWCPP_68 U20 (O[68], I_R[68], S);
  BWCPP_69 U21 (O[69], I_R[69], S);
  BWCPP_70 U22 (O[70], I_R[70], S);
  BWCPP_71 U23 (O[71], I_R[71], S);
  BWCPP_72 U24 (O[72], I_R[72], S);
  BWCPP_73 U25 (O[73], I_R[73], S);
  BWCPP_74 U26 (O[74], I_R[74], S);
  BWCPP_75 U27 (O[75], I_R[75], S);
  BWCPP_76 U28 (O[76], I_R[76], S);
  BWCPP_77 U29 (O[77], I_R[77], S);
  BWCPP_78 U30 (O[78], I_R[78], S);
  BWCPP_79 U31 (O[79], I_R[79], S);
  BWCPP_80 U32 (O[80], I_R[80], S);
  BWCPP_81 U33 (O[81], I_R[81], S);
  BWCPP_82 U34 (O[82], I_R[82], S);
  BWCPP_83 U35 (O[83], I_R[83], S);
  BWCPP_84 U36 (O[84], I_R[84], S);
  BWCPP_85 U37 (O[85], I_R[85], S);
  BWCPP_86 U38 (O[86], I_R[86], S);
  BWCPP_87 U39 (O[87], I_R[87], S);
  BWCPP_88 U40 (O[88], I_R[88], S);
  BWCPP_89 U41 (O[89], I_R[89], S);
  BWCPP_90 U42 (O[90], I_R[90], S);
  BWCPP_91 U43 (O[91], I_R[91], S);
  BWCPP_92 U44 (O[92], I_R[92], S);
  BWCPP_93 U45 (O[93], I_R[93], S);
  BWCPP_94 U46 (O[94], I_R[94], S);
  BWCPP_95 U47 (O[95], I_R[95], S);
  BWCPP_96 U48 (O[96], I_R[96], S);
  BWCPP_97 U49 (O[97], I_R[97], S);
  BWCPP_98 U50 (O[98], I_R[98], S);
  BWCPP_99 U51 (O[99], I_R[99], S);
  BWCPP_100 U52 (O[100], I_R[100], S);
  BWCPP_101 U53 (O[101], I_R[101], S);
  BWCPP_102 U54 (O[102], I_R[102], S);
  BWCPP_103 U55 (O[103], I_R[103], S);
  BWCPP_104 U56 (O[104], I_R[104], S);
  BWCPP_105 U57 (O[105], I_R[105], S);
  BWCPP_106 U58 (O[106], I_R[106], S);
  BWCPP_107 U59 (O[107], I_R[107], S);
  BWCPP_108 U60 (O[108], I_R[108], S);
  BWCPP_109 U61 (O[109], I_R[109], S);
  BWCPP_110 U62 (O[110], I_R[110], S);
  BWCPP_111 U63 (O[111], I_R[111], S);
  BWCNP_112 U64 (O[112], I_T, S);
endmodule

module TUBWCON_114_50 (O, I_T, I_R, S);
  output [114:50] O;
  input [113:50] I_R;
  input I_T;
  input S;
  BWCPP_50 U0 (O[50], I_R[50], S);
  BWCPP_51 U1 (O[51], I_R[51], S);
  BWCPP_52 U2 (O[52], I_R[52], S);
  BWCPP_53 U3 (O[53], I_R[53], S);
  BWCPP_54 U4 (O[54], I_R[54], S);
  BWCPP_55 U5 (O[55], I_R[55], S);
  BWCPP_56 U6 (O[56], I_R[56], S);
  BWCPP_57 U7 (O[57], I_R[57], S);
  BWCPP_58 U8 (O[58], I_R[58], S);
  BWCPP_59 U9 (O[59], I_R[59], S);
  BWCPP_60 U10 (O[60], I_R[60], S);
  BWCPP_61 U11 (O[61], I_R[61], S);
  BWCPP_62 U12 (O[62], I_R[62], S);
  BWCPP_63 U13 (O[63], I_R[63], S);
  BWCPP_64 U14 (O[64], I_R[64], S);
  BWCPP_65 U15 (O[65], I_R[65], S);
  BWCPP_66 U16 (O[66], I_R[66], S);
  BWCPP_67 U17 (O[67], I_R[67], S);
  BWCPP_68 U18 (O[68], I_R[68], S);
  BWCPP_69 U19 (O[69], I_R[69], S);
  BWCPP_70 U20 (O[70], I_R[70], S);
  BWCPP_71 U21 (O[71], I_R[71], S);
  BWCPP_72 U22 (O[72], I_R[72], S);
  BWCPP_73 U23 (O[73], I_R[73], S);
  BWCPP_74 U24 (O[74], I_R[74], S);
  BWCPP_75 U25 (O[75], I_R[75], S);
  BWCPP_76 U26 (O[76], I_R[76], S);
  BWCPP_77 U27 (O[77], I_R[77], S);
  BWCPP_78 U28 (O[78], I_R[78], S);
  BWCPP_79 U29 (O[79], I_R[79], S);
  BWCPP_80 U30 (O[80], I_R[80], S);
  BWCPP_81 U31 (O[81], I_R[81], S);
  BWCPP_82 U32 (O[82], I_R[82], S);
  BWCPP_83 U33 (O[83], I_R[83], S);
  BWCPP_84 U34 (O[84], I_R[84], S);
  BWCPP_85 U35 (O[85], I_R[85], S);
  BWCPP_86 U36 (O[86], I_R[86], S);
  BWCPP_87 U37 (O[87], I_R[87], S);
  BWCPP_88 U38 (O[88], I_R[88], S);
  BWCPP_89 U39 (O[89], I_R[89], S);
  BWCPP_90 U40 (O[90], I_R[90], S);
  BWCPP_91 U41 (O[91], I_R[91], S);
  BWCPP_92 U42 (O[92], I_R[92], S);
  BWCPP_93 U43 (O[93], I_R[93], S);
  BWCPP_94 U44 (O[94], I_R[94], S);
  BWCPP_95 U45 (O[95], I_R[95], S);
  BWCPP_96 U46 (O[96], I_R[96], S);
  BWCPP_97 U47 (O[97], I_R[97], S);
  BWCPP_98 U48 (O[98], I_R[98], S);
  BWCPP_99 U49 (O[99], I_R[99], S);
  BWCPP_100 U50 (O[100], I_R[100], S);
  BWCPP_101 U51 (O[101], I_R[101], S);
  BWCPP_102 U52 (O[102], I_R[102], S);
  BWCPP_103 U53 (O[103], I_R[103], S);
  BWCPP_104 U54 (O[104], I_R[104], S);
  BWCPP_105 U55 (O[105], I_R[105], S);
  BWCPP_106 U56 (O[106], I_R[106], S);
  BWCPP_107 U57 (O[107], I_R[107], S);
  BWCPP_108 U58 (O[108], I_R[108], S);
  BWCPP_109 U59 (O[109], I_R[109], S);
  BWCPP_110 U60 (O[110], I_R[110], S);
  BWCPP_111 U61 (O[111], I_R[111], S);
  BWCPP_112 U62 (O[112], I_R[112], S);
  BWCPP_113 U63 (O[113], I_R[113], S);
  BWCNP_114 U64 (O[114], I_T, S);
endmodule

module TUBWCON_116_52 (O, I_T, I_R, S);
  output [116:52] O;
  input [115:52] I_R;
  input I_T;
  input S;
  BWCPP_52 U0 (O[52], I_R[52], S);
  BWCPP_53 U1 (O[53], I_R[53], S);
  BWCPP_54 U2 (O[54], I_R[54], S);
  BWCPP_55 U3 (O[55], I_R[55], S);
  BWCPP_56 U4 (O[56], I_R[56], S);
  BWCPP_57 U5 (O[57], I_R[57], S);
  BWCPP_58 U6 (O[58], I_R[58], S);
  BWCPP_59 U7 (O[59], I_R[59], S);
  BWCPP_60 U8 (O[60], I_R[60], S);
  BWCPP_61 U9 (O[61], I_R[61], S);
  BWCPP_62 U10 (O[62], I_R[62], S);
  BWCPP_63 U11 (O[63], I_R[63], S);
  BWCPP_64 U12 (O[64], I_R[64], S);
  BWCPP_65 U13 (O[65], I_R[65], S);
  BWCPP_66 U14 (O[66], I_R[66], S);
  BWCPP_67 U15 (O[67], I_R[67], S);
  BWCPP_68 U16 (O[68], I_R[68], S);
  BWCPP_69 U17 (O[69], I_R[69], S);
  BWCPP_70 U18 (O[70], I_R[70], S);
  BWCPP_71 U19 (O[71], I_R[71], S);
  BWCPP_72 U20 (O[72], I_R[72], S);
  BWCPP_73 U21 (O[73], I_R[73], S);
  BWCPP_74 U22 (O[74], I_R[74], S);
  BWCPP_75 U23 (O[75], I_R[75], S);
  BWCPP_76 U24 (O[76], I_R[76], S);
  BWCPP_77 U25 (O[77], I_R[77], S);
  BWCPP_78 U26 (O[78], I_R[78], S);
  BWCPP_79 U27 (O[79], I_R[79], S);
  BWCPP_80 U28 (O[80], I_R[80], S);
  BWCPP_81 U29 (O[81], I_R[81], S);
  BWCPP_82 U30 (O[82], I_R[82], S);
  BWCPP_83 U31 (O[83], I_R[83], S);
  BWCPP_84 U32 (O[84], I_R[84], S);
  BWCPP_85 U33 (O[85], I_R[85], S);
  BWCPP_86 U34 (O[86], I_R[86], S);
  BWCPP_87 U35 (O[87], I_R[87], S);
  BWCPP_88 U36 (O[88], I_R[88], S);
  BWCPP_89 U37 (O[89], I_R[89], S);
  BWCPP_90 U38 (O[90], I_R[90], S);
  BWCPP_91 U39 (O[91], I_R[91], S);
  BWCPP_92 U40 (O[92], I_R[92], S);
  BWCPP_93 U41 (O[93], I_R[93], S);
  BWCPP_94 U42 (O[94], I_R[94], S);
  BWCPP_95 U43 (O[95], I_R[95], S);
  BWCPP_96 U44 (O[96], I_R[96], S);
  BWCPP_97 U45 (O[97], I_R[97], S);
  BWCPP_98 U46 (O[98], I_R[98], S);
  BWCPP_99 U47 (O[99], I_R[99], S);
  BWCPP_100 U48 (O[100], I_R[100], S);
  BWCPP_101 U49 (O[101], I_R[101], S);
  BWCPP_102 U50 (O[102], I_R[102], S);
  BWCPP_103 U51 (O[103], I_R[103], S);
  BWCPP_104 U52 (O[104], I_R[104], S);
  BWCPP_105 U53 (O[105], I_R[105], S);
  BWCPP_106 U54 (O[106], I_R[106], S);
  BWCPP_107 U55 (O[107], I_R[107], S);
  BWCPP_108 U56 (O[108], I_R[108], S);
  BWCPP_109 U57 (O[109], I_R[109], S);
  BWCPP_110 U58 (O[110], I_R[110], S);
  BWCPP_111 U59 (O[111], I_R[111], S);
  BWCPP_112 U60 (O[112], I_R[112], S);
  BWCPP_113 U61 (O[113], I_R[113], S);
  BWCPP_114 U62 (O[114], I_R[114], S);
  BWCPP_115 U63 (O[115], I_R[115], S);
  BWCNP_116 U64 (O[116], I_T, S);
endmodule

module TUBWCON_118_54 (O, I_T, I_R, S);
  output [118:54] O;
  input [117:54] I_R;
  input I_T;
  input S;
  BWCPP_54 U0 (O[54], I_R[54], S);
  BWCPP_55 U1 (O[55], I_R[55], S);
  BWCPP_56 U2 (O[56], I_R[56], S);
  BWCPP_57 U3 (O[57], I_R[57], S);
  BWCPP_58 U4 (O[58], I_R[58], S);
  BWCPP_59 U5 (O[59], I_R[59], S);
  BWCPP_60 U6 (O[60], I_R[60], S);
  BWCPP_61 U7 (O[61], I_R[61], S);
  BWCPP_62 U8 (O[62], I_R[62], S);
  BWCPP_63 U9 (O[63], I_R[63], S);
  BWCPP_64 U10 (O[64], I_R[64], S);
  BWCPP_65 U11 (O[65], I_R[65], S);
  BWCPP_66 U12 (O[66], I_R[66], S);
  BWCPP_67 U13 (O[67], I_R[67], S);
  BWCPP_68 U14 (O[68], I_R[68], S);
  BWCPP_69 U15 (O[69], I_R[69], S);
  BWCPP_70 U16 (O[70], I_R[70], S);
  BWCPP_71 U17 (O[71], I_R[71], S);
  BWCPP_72 U18 (O[72], I_R[72], S);
  BWCPP_73 U19 (O[73], I_R[73], S);
  BWCPP_74 U20 (O[74], I_R[74], S);
  BWCPP_75 U21 (O[75], I_R[75], S);
  BWCPP_76 U22 (O[76], I_R[76], S);
  BWCPP_77 U23 (O[77], I_R[77], S);
  BWCPP_78 U24 (O[78], I_R[78], S);
  BWCPP_79 U25 (O[79], I_R[79], S);
  BWCPP_80 U26 (O[80], I_R[80], S);
  BWCPP_81 U27 (O[81], I_R[81], S);
  BWCPP_82 U28 (O[82], I_R[82], S);
  BWCPP_83 U29 (O[83], I_R[83], S);
  BWCPP_84 U30 (O[84], I_R[84], S);
  BWCPP_85 U31 (O[85], I_R[85], S);
  BWCPP_86 U32 (O[86], I_R[86], S);
  BWCPP_87 U33 (O[87], I_R[87], S);
  BWCPP_88 U34 (O[88], I_R[88], S);
  BWCPP_89 U35 (O[89], I_R[89], S);
  BWCPP_90 U36 (O[90], I_R[90], S);
  BWCPP_91 U37 (O[91], I_R[91], S);
  BWCPP_92 U38 (O[92], I_R[92], S);
  BWCPP_93 U39 (O[93], I_R[93], S);
  BWCPP_94 U40 (O[94], I_R[94], S);
  BWCPP_95 U41 (O[95], I_R[95], S);
  BWCPP_96 U42 (O[96], I_R[96], S);
  BWCPP_97 U43 (O[97], I_R[97], S);
  BWCPP_98 U44 (O[98], I_R[98], S);
  BWCPP_99 U45 (O[99], I_R[99], S);
  BWCPP_100 U46 (O[100], I_R[100], S);
  BWCPP_101 U47 (O[101], I_R[101], S);
  BWCPP_102 U48 (O[102], I_R[102], S);
  BWCPP_103 U49 (O[103], I_R[103], S);
  BWCPP_104 U50 (O[104], I_R[104], S);
  BWCPP_105 U51 (O[105], I_R[105], S);
  BWCPP_106 U52 (O[106], I_R[106], S);
  BWCPP_107 U53 (O[107], I_R[107], S);
  BWCPP_108 U54 (O[108], I_R[108], S);
  BWCPP_109 U55 (O[109], I_R[109], S);
  BWCPP_110 U56 (O[110], I_R[110], S);
  BWCPP_111 U57 (O[111], I_R[111], S);
  BWCPP_112 U58 (O[112], I_R[112], S);
  BWCPP_113 U59 (O[113], I_R[113], S);
  BWCPP_114 U60 (O[114], I_R[114], S);
  BWCPP_115 U61 (O[115], I_R[115], S);
  BWCPP_116 U62 (O[116], I_R[116], S);
  BWCPP_117 U63 (O[117], I_R[117], S);
  BWCNP_118 U64 (O[118], I_T, S);
endmodule

module TUBWCON_120_56 (O, I_T, I_R, S);
  output [120:56] O;
  input [119:56] I_R;
  input I_T;
  input S;
  BWCPP_56 U0 (O[56], I_R[56], S);
  BWCPP_57 U1 (O[57], I_R[57], S);
  BWCPP_58 U2 (O[58], I_R[58], S);
  BWCPP_59 U3 (O[59], I_R[59], S);
  BWCPP_60 U4 (O[60], I_R[60], S);
  BWCPP_61 U5 (O[61], I_R[61], S);
  BWCPP_62 U6 (O[62], I_R[62], S);
  BWCPP_63 U7 (O[63], I_R[63], S);
  BWCPP_64 U8 (O[64], I_R[64], S);
  BWCPP_65 U9 (O[65], I_R[65], S);
  BWCPP_66 U10 (O[66], I_R[66], S);
  BWCPP_67 U11 (O[67], I_R[67], S);
  BWCPP_68 U12 (O[68], I_R[68], S);
  BWCPP_69 U13 (O[69], I_R[69], S);
  BWCPP_70 U14 (O[70], I_R[70], S);
  BWCPP_71 U15 (O[71], I_R[71], S);
  BWCPP_72 U16 (O[72], I_R[72], S);
  BWCPP_73 U17 (O[73], I_R[73], S);
  BWCPP_74 U18 (O[74], I_R[74], S);
  BWCPP_75 U19 (O[75], I_R[75], S);
  BWCPP_76 U20 (O[76], I_R[76], S);
  BWCPP_77 U21 (O[77], I_R[77], S);
  BWCPP_78 U22 (O[78], I_R[78], S);
  BWCPP_79 U23 (O[79], I_R[79], S);
  BWCPP_80 U24 (O[80], I_R[80], S);
  BWCPP_81 U25 (O[81], I_R[81], S);
  BWCPP_82 U26 (O[82], I_R[82], S);
  BWCPP_83 U27 (O[83], I_R[83], S);
  BWCPP_84 U28 (O[84], I_R[84], S);
  BWCPP_85 U29 (O[85], I_R[85], S);
  BWCPP_86 U30 (O[86], I_R[86], S);
  BWCPP_87 U31 (O[87], I_R[87], S);
  BWCPP_88 U32 (O[88], I_R[88], S);
  BWCPP_89 U33 (O[89], I_R[89], S);
  BWCPP_90 U34 (O[90], I_R[90], S);
  BWCPP_91 U35 (O[91], I_R[91], S);
  BWCPP_92 U36 (O[92], I_R[92], S);
  BWCPP_93 U37 (O[93], I_R[93], S);
  BWCPP_94 U38 (O[94], I_R[94], S);
  BWCPP_95 U39 (O[95], I_R[95], S);
  BWCPP_96 U40 (O[96], I_R[96], S);
  BWCPP_97 U41 (O[97], I_R[97], S);
  BWCPP_98 U42 (O[98], I_R[98], S);
  BWCPP_99 U43 (O[99], I_R[99], S);
  BWCPP_100 U44 (O[100], I_R[100], S);
  BWCPP_101 U45 (O[101], I_R[101], S);
  BWCPP_102 U46 (O[102], I_R[102], S);
  BWCPP_103 U47 (O[103], I_R[103], S);
  BWCPP_104 U48 (O[104], I_R[104], S);
  BWCPP_105 U49 (O[105], I_R[105], S);
  BWCPP_106 U50 (O[106], I_R[106], S);
  BWCPP_107 U51 (O[107], I_R[107], S);
  BWCPP_108 U52 (O[108], I_R[108], S);
  BWCPP_109 U53 (O[109], I_R[109], S);
  BWCPP_110 U54 (O[110], I_R[110], S);
  BWCPP_111 U55 (O[111], I_R[111], S);
  BWCPP_112 U56 (O[112], I_R[112], S);
  BWCPP_113 U57 (O[113], I_R[113], S);
  BWCPP_114 U58 (O[114], I_R[114], S);
  BWCPP_115 U59 (O[115], I_R[115], S);
  BWCPP_116 U60 (O[116], I_R[116], S);
  BWCPP_117 U61 (O[117], I_R[117], S);
  BWCPP_118 U62 (O[118], I_R[118], S);
  BWCPP_119 U63 (O[119], I_R[119], S);
  BWCNP_120 U64 (O[120], I_T, S);
endmodule

module TUBWCON_122_58 (O, I_T, I_R, S);
  output [122:58] O;
  input [121:58] I_R;
  input I_T;
  input S;
  BWCPP_58 U0 (O[58], I_R[58], S);
  BWCPP_59 U1 (O[59], I_R[59], S);
  BWCPP_60 U2 (O[60], I_R[60], S);
  BWCPP_61 U3 (O[61], I_R[61], S);
  BWCPP_62 U4 (O[62], I_R[62], S);
  BWCPP_63 U5 (O[63], I_R[63], S);
  BWCPP_64 U6 (O[64], I_R[64], S);
  BWCPP_65 U7 (O[65], I_R[65], S);
  BWCPP_66 U8 (O[66], I_R[66], S);
  BWCPP_67 U9 (O[67], I_R[67], S);
  BWCPP_68 U10 (O[68], I_R[68], S);
  BWCPP_69 U11 (O[69], I_R[69], S);
  BWCPP_70 U12 (O[70], I_R[70], S);
  BWCPP_71 U13 (O[71], I_R[71], S);
  BWCPP_72 U14 (O[72], I_R[72], S);
  BWCPP_73 U15 (O[73], I_R[73], S);
  BWCPP_74 U16 (O[74], I_R[74], S);
  BWCPP_75 U17 (O[75], I_R[75], S);
  BWCPP_76 U18 (O[76], I_R[76], S);
  BWCPP_77 U19 (O[77], I_R[77], S);
  BWCPP_78 U20 (O[78], I_R[78], S);
  BWCPP_79 U21 (O[79], I_R[79], S);
  BWCPP_80 U22 (O[80], I_R[80], S);
  BWCPP_81 U23 (O[81], I_R[81], S);
  BWCPP_82 U24 (O[82], I_R[82], S);
  BWCPP_83 U25 (O[83], I_R[83], S);
  BWCPP_84 U26 (O[84], I_R[84], S);
  BWCPP_85 U27 (O[85], I_R[85], S);
  BWCPP_86 U28 (O[86], I_R[86], S);
  BWCPP_87 U29 (O[87], I_R[87], S);
  BWCPP_88 U30 (O[88], I_R[88], S);
  BWCPP_89 U31 (O[89], I_R[89], S);
  BWCPP_90 U32 (O[90], I_R[90], S);
  BWCPP_91 U33 (O[91], I_R[91], S);
  BWCPP_92 U34 (O[92], I_R[92], S);
  BWCPP_93 U35 (O[93], I_R[93], S);
  BWCPP_94 U36 (O[94], I_R[94], S);
  BWCPP_95 U37 (O[95], I_R[95], S);
  BWCPP_96 U38 (O[96], I_R[96], S);
  BWCPP_97 U39 (O[97], I_R[97], S);
  BWCPP_98 U40 (O[98], I_R[98], S);
  BWCPP_99 U41 (O[99], I_R[99], S);
  BWCPP_100 U42 (O[100], I_R[100], S);
  BWCPP_101 U43 (O[101], I_R[101], S);
  BWCPP_102 U44 (O[102], I_R[102], S);
  BWCPP_103 U45 (O[103], I_R[103], S);
  BWCPP_104 U46 (O[104], I_R[104], S);
  BWCPP_105 U47 (O[105], I_R[105], S);
  BWCPP_106 U48 (O[106], I_R[106], S);
  BWCPP_107 U49 (O[107], I_R[107], S);
  BWCPP_108 U50 (O[108], I_R[108], S);
  BWCPP_109 U51 (O[109], I_R[109], S);
  BWCPP_110 U52 (O[110], I_R[110], S);
  BWCPP_111 U53 (O[111], I_R[111], S);
  BWCPP_112 U54 (O[112], I_R[112], S);
  BWCPP_113 U55 (O[113], I_R[113], S);
  BWCPP_114 U56 (O[114], I_R[114], S);
  BWCPP_115 U57 (O[115], I_R[115], S);
  BWCPP_116 U58 (O[116], I_R[116], S);
  BWCPP_117 U59 (O[117], I_R[117], S);
  BWCPP_118 U60 (O[118], I_R[118], S);
  BWCPP_119 U61 (O[119], I_R[119], S);
  BWCPP_120 U62 (O[120], I_R[120], S);
  BWCPP_121 U63 (O[121], I_R[121], S);
  BWCNP_122 U64 (O[122], I_T, S);
endmodule

module TUBWCON_124_60 (O, I_T, I_R, S);
  output [124:60] O;
  input [123:60] I_R;
  input I_T;
  input S;
  BWCPP_60 U0 (O[60], I_R[60], S);
  BWCPP_61 U1 (O[61], I_R[61], S);
  BWCPP_62 U2 (O[62], I_R[62], S);
  BWCPP_63 U3 (O[63], I_R[63], S);
  BWCPP_64 U4 (O[64], I_R[64], S);
  BWCPP_65 U5 (O[65], I_R[65], S);
  BWCPP_66 U6 (O[66], I_R[66], S);
  BWCPP_67 U7 (O[67], I_R[67], S);
  BWCPP_68 U8 (O[68], I_R[68], S);
  BWCPP_69 U9 (O[69], I_R[69], S);
  BWCPP_70 U10 (O[70], I_R[70], S);
  BWCPP_71 U11 (O[71], I_R[71], S);
  BWCPP_72 U12 (O[72], I_R[72], S);
  BWCPP_73 U13 (O[73], I_R[73], S);
  BWCPP_74 U14 (O[74], I_R[74], S);
  BWCPP_75 U15 (O[75], I_R[75], S);
  BWCPP_76 U16 (O[76], I_R[76], S);
  BWCPP_77 U17 (O[77], I_R[77], S);
  BWCPP_78 U18 (O[78], I_R[78], S);
  BWCPP_79 U19 (O[79], I_R[79], S);
  BWCPP_80 U20 (O[80], I_R[80], S);
  BWCPP_81 U21 (O[81], I_R[81], S);
  BWCPP_82 U22 (O[82], I_R[82], S);
  BWCPP_83 U23 (O[83], I_R[83], S);
  BWCPP_84 U24 (O[84], I_R[84], S);
  BWCPP_85 U25 (O[85], I_R[85], S);
  BWCPP_86 U26 (O[86], I_R[86], S);
  BWCPP_87 U27 (O[87], I_R[87], S);
  BWCPP_88 U28 (O[88], I_R[88], S);
  BWCPP_89 U29 (O[89], I_R[89], S);
  BWCPP_90 U30 (O[90], I_R[90], S);
  BWCPP_91 U31 (O[91], I_R[91], S);
  BWCPP_92 U32 (O[92], I_R[92], S);
  BWCPP_93 U33 (O[93], I_R[93], S);
  BWCPP_94 U34 (O[94], I_R[94], S);
  BWCPP_95 U35 (O[95], I_R[95], S);
  BWCPP_96 U36 (O[96], I_R[96], S);
  BWCPP_97 U37 (O[97], I_R[97], S);
  BWCPP_98 U38 (O[98], I_R[98], S);
  BWCPP_99 U39 (O[99], I_R[99], S);
  BWCPP_100 U40 (O[100], I_R[100], S);
  BWCPP_101 U41 (O[101], I_R[101], S);
  BWCPP_102 U42 (O[102], I_R[102], S);
  BWCPP_103 U43 (O[103], I_R[103], S);
  BWCPP_104 U44 (O[104], I_R[104], S);
  BWCPP_105 U45 (O[105], I_R[105], S);
  BWCPP_106 U46 (O[106], I_R[106], S);
  BWCPP_107 U47 (O[107], I_R[107], S);
  BWCPP_108 U48 (O[108], I_R[108], S);
  BWCPP_109 U49 (O[109], I_R[109], S);
  BWCPP_110 U50 (O[110], I_R[110], S);
  BWCPP_111 U51 (O[111], I_R[111], S);
  BWCPP_112 U52 (O[112], I_R[112], S);
  BWCPP_113 U53 (O[113], I_R[113], S);
  BWCPP_114 U54 (O[114], I_R[114], S);
  BWCPP_115 U55 (O[115], I_R[115], S);
  BWCPP_116 U56 (O[116], I_R[116], S);
  BWCPP_117 U57 (O[117], I_R[117], S);
  BWCPP_118 U58 (O[118], I_R[118], S);
  BWCPP_119 U59 (O[119], I_R[119], S);
  BWCPP_120 U60 (O[120], I_R[120], S);
  BWCPP_121 U61 (O[121], I_R[121], S);
  BWCPP_122 U62 (O[122], I_R[122], S);
  BWCPP_123 U63 (O[123], I_R[123], S);
  BWCNP_124 U64 (O[124], I_T, S);
endmodule

module TUBWCON_126_62 (O, I_T, I_R, S);
  output [126:62] O;
  input [125:62] I_R;
  input I_T;
  input S;
  BWCPP_62 U0 (O[62], I_R[62], S);
  BWCPP_63 U1 (O[63], I_R[63], S);
  BWCPP_64 U2 (O[64], I_R[64], S);
  BWCPP_65 U3 (O[65], I_R[65], S);
  BWCPP_66 U4 (O[66], I_R[66], S);
  BWCPP_67 U5 (O[67], I_R[67], S);
  BWCPP_68 U6 (O[68], I_R[68], S);
  BWCPP_69 U7 (O[69], I_R[69], S);
  BWCPP_70 U8 (O[70], I_R[70], S);
  BWCPP_71 U9 (O[71], I_R[71], S);
  BWCPP_72 U10 (O[72], I_R[72], S);
  BWCPP_73 U11 (O[73], I_R[73], S);
  BWCPP_74 U12 (O[74], I_R[74], S);
  BWCPP_75 U13 (O[75], I_R[75], S);
  BWCPP_76 U14 (O[76], I_R[76], S);
  BWCPP_77 U15 (O[77], I_R[77], S);
  BWCPP_78 U16 (O[78], I_R[78], S);
  BWCPP_79 U17 (O[79], I_R[79], S);
  BWCPP_80 U18 (O[80], I_R[80], S);
  BWCPP_81 U19 (O[81], I_R[81], S);
  BWCPP_82 U20 (O[82], I_R[82], S);
  BWCPP_83 U21 (O[83], I_R[83], S);
  BWCPP_84 U22 (O[84], I_R[84], S);
  BWCPP_85 U23 (O[85], I_R[85], S);
  BWCPP_86 U24 (O[86], I_R[86], S);
  BWCPP_87 U25 (O[87], I_R[87], S);
  BWCPP_88 U26 (O[88], I_R[88], S);
  BWCPP_89 U27 (O[89], I_R[89], S);
  BWCPP_90 U28 (O[90], I_R[90], S);
  BWCPP_91 U29 (O[91], I_R[91], S);
  BWCPP_92 U30 (O[92], I_R[92], S);
  BWCPP_93 U31 (O[93], I_R[93], S);
  BWCPP_94 U32 (O[94], I_R[94], S);
  BWCPP_95 U33 (O[95], I_R[95], S);
  BWCPP_96 U34 (O[96], I_R[96], S);
  BWCPP_97 U35 (O[97], I_R[97], S);
  BWCPP_98 U36 (O[98], I_R[98], S);
  BWCPP_99 U37 (O[99], I_R[99], S);
  BWCPP_100 U38 (O[100], I_R[100], S);
  BWCPP_101 U39 (O[101], I_R[101], S);
  BWCPP_102 U40 (O[102], I_R[102], S);
  BWCPP_103 U41 (O[103], I_R[103], S);
  BWCPP_104 U42 (O[104], I_R[104], S);
  BWCPP_105 U43 (O[105], I_R[105], S);
  BWCPP_106 U44 (O[106], I_R[106], S);
  BWCPP_107 U45 (O[107], I_R[107], S);
  BWCPP_108 U46 (O[108], I_R[108], S);
  BWCPP_109 U47 (O[109], I_R[109], S);
  BWCPP_110 U48 (O[110], I_R[110], S);
  BWCPP_111 U49 (O[111], I_R[111], S);
  BWCPP_112 U50 (O[112], I_R[112], S);
  BWCPP_113 U51 (O[113], I_R[113], S);
  BWCPP_114 U52 (O[114], I_R[114], S);
  BWCPP_115 U53 (O[115], I_R[115], S);
  BWCPP_116 U54 (O[116], I_R[116], S);
  BWCPP_117 U55 (O[117], I_R[117], S);
  BWCPP_118 U56 (O[118], I_R[118], S);
  BWCPP_119 U57 (O[119], I_R[119], S);
  BWCPP_120 U58 (O[120], I_R[120], S);
  BWCPP_121 U59 (O[121], I_R[121], S);
  BWCPP_122 U60 (O[122], I_R[122], S);
  BWCPP_123 U61 (O[123], I_R[123], S);
  BWCPP_124 U62 (O[124], I_R[124], S);
  BWCPP_125 U63 (O[125], I_R[125], S);
  BWCNP_126 U64 (O[126], I_T, S);
endmodule

module TUBWCON_64_0 (O, I_T, I_R, S);
  output [64:0] O;
  input [63:0] I_R;
  input I_T;
  input S;
  BWCPP_0 U0 (O[0], I_R[0], S);
  BWCPP_1 U1 (O[1], I_R[1], S);
  BWCPP_2 U2 (O[2], I_R[2], S);
  BWCPP_3 U3 (O[3], I_R[3], S);
  BWCPP_4 U4 (O[4], I_R[4], S);
  BWCPP_5 U5 (O[5], I_R[5], S);
  BWCPP_6 U6 (O[6], I_R[6], S);
  BWCPP_7 U7 (O[7], I_R[7], S);
  BWCPP_8 U8 (O[8], I_R[8], S);
  BWCPP_9 U9 (O[9], I_R[9], S);
  BWCPP_10 U10 (O[10], I_R[10], S);
  BWCPP_11 U11 (O[11], I_R[11], S);
  BWCPP_12 U12 (O[12], I_R[12], S);
  BWCPP_13 U13 (O[13], I_R[13], S);
  BWCPP_14 U14 (O[14], I_R[14], S);
  BWCPP_15 U15 (O[15], I_R[15], S);
  BWCPP_16 U16 (O[16], I_R[16], S);
  BWCPP_17 U17 (O[17], I_R[17], S);
  BWCPP_18 U18 (O[18], I_R[18], S);
  BWCPP_19 U19 (O[19], I_R[19], S);
  BWCPP_20 U20 (O[20], I_R[20], S);
  BWCPP_21 U21 (O[21], I_R[21], S);
  BWCPP_22 U22 (O[22], I_R[22], S);
  BWCPP_23 U23 (O[23], I_R[23], S);
  BWCPP_24 U24 (O[24], I_R[24], S);
  BWCPP_25 U25 (O[25], I_R[25], S);
  BWCPP_26 U26 (O[26], I_R[26], S);
  BWCPP_27 U27 (O[27], I_R[27], S);
  BWCPP_28 U28 (O[28], I_R[28], S);
  BWCPP_29 U29 (O[29], I_R[29], S);
  BWCPP_30 U30 (O[30], I_R[30], S);
  BWCPP_31 U31 (O[31], I_R[31], S);
  BWCPP_32 U32 (O[32], I_R[32], S);
  BWCPP_33 U33 (O[33], I_R[33], S);
  BWCPP_34 U34 (O[34], I_R[34], S);
  BWCPP_35 U35 (O[35], I_R[35], S);
  BWCPP_36 U36 (O[36], I_R[36], S);
  BWCPP_37 U37 (O[37], I_R[37], S);
  BWCPP_38 U38 (O[38], I_R[38], S);
  BWCPP_39 U39 (O[39], I_R[39], S);
  BWCPP_40 U40 (O[40], I_R[40], S);
  BWCPP_41 U41 (O[41], I_R[41], S);
  BWCPP_42 U42 (O[42], I_R[42], S);
  BWCPP_43 U43 (O[43], I_R[43], S);
  BWCPP_44 U44 (O[44], I_R[44], S);
  BWCPP_45 U45 (O[45], I_R[45], S);
  BWCPP_46 U46 (O[46], I_R[46], S);
  BWCPP_47 U47 (O[47], I_R[47], S);
  BWCPP_48 U48 (O[48], I_R[48], S);
  BWCPP_49 U49 (O[49], I_R[49], S);
  BWCPP_50 U50 (O[50], I_R[50], S);
  BWCPP_51 U51 (O[51], I_R[51], S);
  BWCPP_52 U52 (O[52], I_R[52], S);
  BWCPP_53 U53 (O[53], I_R[53], S);
  BWCPP_54 U54 (O[54], I_R[54], S);
  BWCPP_55 U55 (O[55], I_R[55], S);
  BWCPP_56 U56 (O[56], I_R[56], S);
  BWCPP_57 U57 (O[57], I_R[57], S);
  BWCPP_58 U58 (O[58], I_R[58], S);
  BWCPP_59 U59 (O[59], I_R[59], S);
  BWCPP_60 U60 (O[60], I_R[60], S);
  BWCPP_61 U61 (O[61], I_R[61], S);
  BWCPP_62 U62 (O[62], I_R[62], S);
  BWCPP_63 U63 (O[63], I_R[63], S);
  BWCNP_64 U64 (O[64], I_T, S);
endmodule

module TUBWCON_66_2 (O, I_T, I_R, S);
  output [66:2] O;
  input [65:2] I_R;
  input I_T;
  input S;
  BWCPP_2 U0 (O[2], I_R[2], S);
  BWCPP_3 U1 (O[3], I_R[3], S);
  BWCPP_4 U2 (O[4], I_R[4], S);
  BWCPP_5 U3 (O[5], I_R[5], S);
  BWCPP_6 U4 (O[6], I_R[6], S);
  BWCPP_7 U5 (O[7], I_R[7], S);
  BWCPP_8 U6 (O[8], I_R[8], S);
  BWCPP_9 U7 (O[9], I_R[9], S);
  BWCPP_10 U8 (O[10], I_R[10], S);
  BWCPP_11 U9 (O[11], I_R[11], S);
  BWCPP_12 U10 (O[12], I_R[12], S);
  BWCPP_13 U11 (O[13], I_R[13], S);
  BWCPP_14 U12 (O[14], I_R[14], S);
  BWCPP_15 U13 (O[15], I_R[15], S);
  BWCPP_16 U14 (O[16], I_R[16], S);
  BWCPP_17 U15 (O[17], I_R[17], S);
  BWCPP_18 U16 (O[18], I_R[18], S);
  BWCPP_19 U17 (O[19], I_R[19], S);
  BWCPP_20 U18 (O[20], I_R[20], S);
  BWCPP_21 U19 (O[21], I_R[21], S);
  BWCPP_22 U20 (O[22], I_R[22], S);
  BWCPP_23 U21 (O[23], I_R[23], S);
  BWCPP_24 U22 (O[24], I_R[24], S);
  BWCPP_25 U23 (O[25], I_R[25], S);
  BWCPP_26 U24 (O[26], I_R[26], S);
  BWCPP_27 U25 (O[27], I_R[27], S);
  BWCPP_28 U26 (O[28], I_R[28], S);
  BWCPP_29 U27 (O[29], I_R[29], S);
  BWCPP_30 U28 (O[30], I_R[30], S);
  BWCPP_31 U29 (O[31], I_R[31], S);
  BWCPP_32 U30 (O[32], I_R[32], S);
  BWCPP_33 U31 (O[33], I_R[33], S);
  BWCPP_34 U32 (O[34], I_R[34], S);
  BWCPP_35 U33 (O[35], I_R[35], S);
  BWCPP_36 U34 (O[36], I_R[36], S);
  BWCPP_37 U35 (O[37], I_R[37], S);
  BWCPP_38 U36 (O[38], I_R[38], S);
  BWCPP_39 U37 (O[39], I_R[39], S);
  BWCPP_40 U38 (O[40], I_R[40], S);
  BWCPP_41 U39 (O[41], I_R[41], S);
  BWCPP_42 U40 (O[42], I_R[42], S);
  BWCPP_43 U41 (O[43], I_R[43], S);
  BWCPP_44 U42 (O[44], I_R[44], S);
  BWCPP_45 U43 (O[45], I_R[45], S);
  BWCPP_46 U44 (O[46], I_R[46], S);
  BWCPP_47 U45 (O[47], I_R[47], S);
  BWCPP_48 U46 (O[48], I_R[48], S);
  BWCPP_49 U47 (O[49], I_R[49], S);
  BWCPP_50 U48 (O[50], I_R[50], S);
  BWCPP_51 U49 (O[51], I_R[51], S);
  BWCPP_52 U50 (O[52], I_R[52], S);
  BWCPP_53 U51 (O[53], I_R[53], S);
  BWCPP_54 U52 (O[54], I_R[54], S);
  BWCPP_55 U53 (O[55], I_R[55], S);
  BWCPP_56 U54 (O[56], I_R[56], S);
  BWCPP_57 U55 (O[57], I_R[57], S);
  BWCPP_58 U56 (O[58], I_R[58], S);
  BWCPP_59 U57 (O[59], I_R[59], S);
  BWCPP_60 U58 (O[60], I_R[60], S);
  BWCPP_61 U59 (O[61], I_R[61], S);
  BWCPP_62 U60 (O[62], I_R[62], S);
  BWCPP_63 U61 (O[63], I_R[63], S);
  BWCPP_64 U62 (O[64], I_R[64], S);
  BWCPP_65 U63 (O[65], I_R[65], S);
  BWCNP_66 U64 (O[66], I_T, S);
endmodule

module TUBWCON_68_4 (O, I_T, I_R, S);
  output [68:4] O;
  input [67:4] I_R;
  input I_T;
  input S;
  BWCPP_4 U0 (O[4], I_R[4], S);
  BWCPP_5 U1 (O[5], I_R[5], S);
  BWCPP_6 U2 (O[6], I_R[6], S);
  BWCPP_7 U3 (O[7], I_R[7], S);
  BWCPP_8 U4 (O[8], I_R[8], S);
  BWCPP_9 U5 (O[9], I_R[9], S);
  BWCPP_10 U6 (O[10], I_R[10], S);
  BWCPP_11 U7 (O[11], I_R[11], S);
  BWCPP_12 U8 (O[12], I_R[12], S);
  BWCPP_13 U9 (O[13], I_R[13], S);
  BWCPP_14 U10 (O[14], I_R[14], S);
  BWCPP_15 U11 (O[15], I_R[15], S);
  BWCPP_16 U12 (O[16], I_R[16], S);
  BWCPP_17 U13 (O[17], I_R[17], S);
  BWCPP_18 U14 (O[18], I_R[18], S);
  BWCPP_19 U15 (O[19], I_R[19], S);
  BWCPP_20 U16 (O[20], I_R[20], S);
  BWCPP_21 U17 (O[21], I_R[21], S);
  BWCPP_22 U18 (O[22], I_R[22], S);
  BWCPP_23 U19 (O[23], I_R[23], S);
  BWCPP_24 U20 (O[24], I_R[24], S);
  BWCPP_25 U21 (O[25], I_R[25], S);
  BWCPP_26 U22 (O[26], I_R[26], S);
  BWCPP_27 U23 (O[27], I_R[27], S);
  BWCPP_28 U24 (O[28], I_R[28], S);
  BWCPP_29 U25 (O[29], I_R[29], S);
  BWCPP_30 U26 (O[30], I_R[30], S);
  BWCPP_31 U27 (O[31], I_R[31], S);
  BWCPP_32 U28 (O[32], I_R[32], S);
  BWCPP_33 U29 (O[33], I_R[33], S);
  BWCPP_34 U30 (O[34], I_R[34], S);
  BWCPP_35 U31 (O[35], I_R[35], S);
  BWCPP_36 U32 (O[36], I_R[36], S);
  BWCPP_37 U33 (O[37], I_R[37], S);
  BWCPP_38 U34 (O[38], I_R[38], S);
  BWCPP_39 U35 (O[39], I_R[39], S);
  BWCPP_40 U36 (O[40], I_R[40], S);
  BWCPP_41 U37 (O[41], I_R[41], S);
  BWCPP_42 U38 (O[42], I_R[42], S);
  BWCPP_43 U39 (O[43], I_R[43], S);
  BWCPP_44 U40 (O[44], I_R[44], S);
  BWCPP_45 U41 (O[45], I_R[45], S);
  BWCPP_46 U42 (O[46], I_R[46], S);
  BWCPP_47 U43 (O[47], I_R[47], S);
  BWCPP_48 U44 (O[48], I_R[48], S);
  BWCPP_49 U45 (O[49], I_R[49], S);
  BWCPP_50 U46 (O[50], I_R[50], S);
  BWCPP_51 U47 (O[51], I_R[51], S);
  BWCPP_52 U48 (O[52], I_R[52], S);
  BWCPP_53 U49 (O[53], I_R[53], S);
  BWCPP_54 U50 (O[54], I_R[54], S);
  BWCPP_55 U51 (O[55], I_R[55], S);
  BWCPP_56 U52 (O[56], I_R[56], S);
  BWCPP_57 U53 (O[57], I_R[57], S);
  BWCPP_58 U54 (O[58], I_R[58], S);
  BWCPP_59 U55 (O[59], I_R[59], S);
  BWCPP_60 U56 (O[60], I_R[60], S);
  BWCPP_61 U57 (O[61], I_R[61], S);
  BWCPP_62 U58 (O[62], I_R[62], S);
  BWCPP_63 U59 (O[63], I_R[63], S);
  BWCPP_64 U60 (O[64], I_R[64], S);
  BWCPP_65 U61 (O[65], I_R[65], S);
  BWCPP_66 U62 (O[66], I_R[66], S);
  BWCPP_67 U63 (O[67], I_R[67], S);
  BWCNP_68 U64 (O[68], I_T, S);
endmodule

module TUBWCON_70_6 (O, I_T, I_R, S);
  output [70:6] O;
  input [69:6] I_R;
  input I_T;
  input S;
  BWCPP_6 U0 (O[6], I_R[6], S);
  BWCPP_7 U1 (O[7], I_R[7], S);
  BWCPP_8 U2 (O[8], I_R[8], S);
  BWCPP_9 U3 (O[9], I_R[9], S);
  BWCPP_10 U4 (O[10], I_R[10], S);
  BWCPP_11 U5 (O[11], I_R[11], S);
  BWCPP_12 U6 (O[12], I_R[12], S);
  BWCPP_13 U7 (O[13], I_R[13], S);
  BWCPP_14 U8 (O[14], I_R[14], S);
  BWCPP_15 U9 (O[15], I_R[15], S);
  BWCPP_16 U10 (O[16], I_R[16], S);
  BWCPP_17 U11 (O[17], I_R[17], S);
  BWCPP_18 U12 (O[18], I_R[18], S);
  BWCPP_19 U13 (O[19], I_R[19], S);
  BWCPP_20 U14 (O[20], I_R[20], S);
  BWCPP_21 U15 (O[21], I_R[21], S);
  BWCPP_22 U16 (O[22], I_R[22], S);
  BWCPP_23 U17 (O[23], I_R[23], S);
  BWCPP_24 U18 (O[24], I_R[24], S);
  BWCPP_25 U19 (O[25], I_R[25], S);
  BWCPP_26 U20 (O[26], I_R[26], S);
  BWCPP_27 U21 (O[27], I_R[27], S);
  BWCPP_28 U22 (O[28], I_R[28], S);
  BWCPP_29 U23 (O[29], I_R[29], S);
  BWCPP_30 U24 (O[30], I_R[30], S);
  BWCPP_31 U25 (O[31], I_R[31], S);
  BWCPP_32 U26 (O[32], I_R[32], S);
  BWCPP_33 U27 (O[33], I_R[33], S);
  BWCPP_34 U28 (O[34], I_R[34], S);
  BWCPP_35 U29 (O[35], I_R[35], S);
  BWCPP_36 U30 (O[36], I_R[36], S);
  BWCPP_37 U31 (O[37], I_R[37], S);
  BWCPP_38 U32 (O[38], I_R[38], S);
  BWCPP_39 U33 (O[39], I_R[39], S);
  BWCPP_40 U34 (O[40], I_R[40], S);
  BWCPP_41 U35 (O[41], I_R[41], S);
  BWCPP_42 U36 (O[42], I_R[42], S);
  BWCPP_43 U37 (O[43], I_R[43], S);
  BWCPP_44 U38 (O[44], I_R[44], S);
  BWCPP_45 U39 (O[45], I_R[45], S);
  BWCPP_46 U40 (O[46], I_R[46], S);
  BWCPP_47 U41 (O[47], I_R[47], S);
  BWCPP_48 U42 (O[48], I_R[48], S);
  BWCPP_49 U43 (O[49], I_R[49], S);
  BWCPP_50 U44 (O[50], I_R[50], S);
  BWCPP_51 U45 (O[51], I_R[51], S);
  BWCPP_52 U46 (O[52], I_R[52], S);
  BWCPP_53 U47 (O[53], I_R[53], S);
  BWCPP_54 U48 (O[54], I_R[54], S);
  BWCPP_55 U49 (O[55], I_R[55], S);
  BWCPP_56 U50 (O[56], I_R[56], S);
  BWCPP_57 U51 (O[57], I_R[57], S);
  BWCPP_58 U52 (O[58], I_R[58], S);
  BWCPP_59 U53 (O[59], I_R[59], S);
  BWCPP_60 U54 (O[60], I_R[60], S);
  BWCPP_61 U55 (O[61], I_R[61], S);
  BWCPP_62 U56 (O[62], I_R[62], S);
  BWCPP_63 U57 (O[63], I_R[63], S);
  BWCPP_64 U58 (O[64], I_R[64], S);
  BWCPP_65 U59 (O[65], I_R[65], S);
  BWCPP_66 U60 (O[66], I_R[66], S);
  BWCPP_67 U61 (O[67], I_R[67], S);
  BWCPP_68 U62 (O[68], I_R[68], S);
  BWCPP_69 U63 (O[69], I_R[69], S);
  BWCNP_70 U64 (O[70], I_T, S);
endmodule

module TUBWCON_72_8 (O, I_T, I_R, S);
  output [72:8] O;
  input [71:8] I_R;
  input I_T;
  input S;
  BWCPP_8 U0 (O[8], I_R[8], S);
  BWCPP_9 U1 (O[9], I_R[9], S);
  BWCPP_10 U2 (O[10], I_R[10], S);
  BWCPP_11 U3 (O[11], I_R[11], S);
  BWCPP_12 U4 (O[12], I_R[12], S);
  BWCPP_13 U5 (O[13], I_R[13], S);
  BWCPP_14 U6 (O[14], I_R[14], S);
  BWCPP_15 U7 (O[15], I_R[15], S);
  BWCPP_16 U8 (O[16], I_R[16], S);
  BWCPP_17 U9 (O[17], I_R[17], S);
  BWCPP_18 U10 (O[18], I_R[18], S);
  BWCPP_19 U11 (O[19], I_R[19], S);
  BWCPP_20 U12 (O[20], I_R[20], S);
  BWCPP_21 U13 (O[21], I_R[21], S);
  BWCPP_22 U14 (O[22], I_R[22], S);
  BWCPP_23 U15 (O[23], I_R[23], S);
  BWCPP_24 U16 (O[24], I_R[24], S);
  BWCPP_25 U17 (O[25], I_R[25], S);
  BWCPP_26 U18 (O[26], I_R[26], S);
  BWCPP_27 U19 (O[27], I_R[27], S);
  BWCPP_28 U20 (O[28], I_R[28], S);
  BWCPP_29 U21 (O[29], I_R[29], S);
  BWCPP_30 U22 (O[30], I_R[30], S);
  BWCPP_31 U23 (O[31], I_R[31], S);
  BWCPP_32 U24 (O[32], I_R[32], S);
  BWCPP_33 U25 (O[33], I_R[33], S);
  BWCPP_34 U26 (O[34], I_R[34], S);
  BWCPP_35 U27 (O[35], I_R[35], S);
  BWCPP_36 U28 (O[36], I_R[36], S);
  BWCPP_37 U29 (O[37], I_R[37], S);
  BWCPP_38 U30 (O[38], I_R[38], S);
  BWCPP_39 U31 (O[39], I_R[39], S);
  BWCPP_40 U32 (O[40], I_R[40], S);
  BWCPP_41 U33 (O[41], I_R[41], S);
  BWCPP_42 U34 (O[42], I_R[42], S);
  BWCPP_43 U35 (O[43], I_R[43], S);
  BWCPP_44 U36 (O[44], I_R[44], S);
  BWCPP_45 U37 (O[45], I_R[45], S);
  BWCPP_46 U38 (O[46], I_R[46], S);
  BWCPP_47 U39 (O[47], I_R[47], S);
  BWCPP_48 U40 (O[48], I_R[48], S);
  BWCPP_49 U41 (O[49], I_R[49], S);
  BWCPP_50 U42 (O[50], I_R[50], S);
  BWCPP_51 U43 (O[51], I_R[51], S);
  BWCPP_52 U44 (O[52], I_R[52], S);
  BWCPP_53 U45 (O[53], I_R[53], S);
  BWCPP_54 U46 (O[54], I_R[54], S);
  BWCPP_55 U47 (O[55], I_R[55], S);
  BWCPP_56 U48 (O[56], I_R[56], S);
  BWCPP_57 U49 (O[57], I_R[57], S);
  BWCPP_58 U50 (O[58], I_R[58], S);
  BWCPP_59 U51 (O[59], I_R[59], S);
  BWCPP_60 U52 (O[60], I_R[60], S);
  BWCPP_61 U53 (O[61], I_R[61], S);
  BWCPP_62 U54 (O[62], I_R[62], S);
  BWCPP_63 U55 (O[63], I_R[63], S);
  BWCPP_64 U56 (O[64], I_R[64], S);
  BWCPP_65 U57 (O[65], I_R[65], S);
  BWCPP_66 U58 (O[66], I_R[66], S);
  BWCPP_67 U59 (O[67], I_R[67], S);
  BWCPP_68 U60 (O[68], I_R[68], S);
  BWCPP_69 U61 (O[69], I_R[69], S);
  BWCPP_70 U62 (O[70], I_R[70], S);
  BWCPP_71 U63 (O[71], I_R[71], S);
  BWCNP_72 U64 (O[72], I_T, S);
endmodule

module TUBWCON_74_10 (O, I_T, I_R, S);
  output [74:10] O;
  input [73:10] I_R;
  input I_T;
  input S;
  BWCPP_10 U0 (O[10], I_R[10], S);
  BWCPP_11 U1 (O[11], I_R[11], S);
  BWCPP_12 U2 (O[12], I_R[12], S);
  BWCPP_13 U3 (O[13], I_R[13], S);
  BWCPP_14 U4 (O[14], I_R[14], S);
  BWCPP_15 U5 (O[15], I_R[15], S);
  BWCPP_16 U6 (O[16], I_R[16], S);
  BWCPP_17 U7 (O[17], I_R[17], S);
  BWCPP_18 U8 (O[18], I_R[18], S);
  BWCPP_19 U9 (O[19], I_R[19], S);
  BWCPP_20 U10 (O[20], I_R[20], S);
  BWCPP_21 U11 (O[21], I_R[21], S);
  BWCPP_22 U12 (O[22], I_R[22], S);
  BWCPP_23 U13 (O[23], I_R[23], S);
  BWCPP_24 U14 (O[24], I_R[24], S);
  BWCPP_25 U15 (O[25], I_R[25], S);
  BWCPP_26 U16 (O[26], I_R[26], S);
  BWCPP_27 U17 (O[27], I_R[27], S);
  BWCPP_28 U18 (O[28], I_R[28], S);
  BWCPP_29 U19 (O[29], I_R[29], S);
  BWCPP_30 U20 (O[30], I_R[30], S);
  BWCPP_31 U21 (O[31], I_R[31], S);
  BWCPP_32 U22 (O[32], I_R[32], S);
  BWCPP_33 U23 (O[33], I_R[33], S);
  BWCPP_34 U24 (O[34], I_R[34], S);
  BWCPP_35 U25 (O[35], I_R[35], S);
  BWCPP_36 U26 (O[36], I_R[36], S);
  BWCPP_37 U27 (O[37], I_R[37], S);
  BWCPP_38 U28 (O[38], I_R[38], S);
  BWCPP_39 U29 (O[39], I_R[39], S);
  BWCPP_40 U30 (O[40], I_R[40], S);
  BWCPP_41 U31 (O[41], I_R[41], S);
  BWCPP_42 U32 (O[42], I_R[42], S);
  BWCPP_43 U33 (O[43], I_R[43], S);
  BWCPP_44 U34 (O[44], I_R[44], S);
  BWCPP_45 U35 (O[45], I_R[45], S);
  BWCPP_46 U36 (O[46], I_R[46], S);
  BWCPP_47 U37 (O[47], I_R[47], S);
  BWCPP_48 U38 (O[48], I_R[48], S);
  BWCPP_49 U39 (O[49], I_R[49], S);
  BWCPP_50 U40 (O[50], I_R[50], S);
  BWCPP_51 U41 (O[51], I_R[51], S);
  BWCPP_52 U42 (O[52], I_R[52], S);
  BWCPP_53 U43 (O[53], I_R[53], S);
  BWCPP_54 U44 (O[54], I_R[54], S);
  BWCPP_55 U45 (O[55], I_R[55], S);
  BWCPP_56 U46 (O[56], I_R[56], S);
  BWCPP_57 U47 (O[57], I_R[57], S);
  BWCPP_58 U48 (O[58], I_R[58], S);
  BWCPP_59 U49 (O[59], I_R[59], S);
  BWCPP_60 U50 (O[60], I_R[60], S);
  BWCPP_61 U51 (O[61], I_R[61], S);
  BWCPP_62 U52 (O[62], I_R[62], S);
  BWCPP_63 U53 (O[63], I_R[63], S);
  BWCPP_64 U54 (O[64], I_R[64], S);
  BWCPP_65 U55 (O[65], I_R[65], S);
  BWCPP_66 U56 (O[66], I_R[66], S);
  BWCPP_67 U57 (O[67], I_R[67], S);
  BWCPP_68 U58 (O[68], I_R[68], S);
  BWCPP_69 U59 (O[69], I_R[69], S);
  BWCPP_70 U60 (O[70], I_R[70], S);
  BWCPP_71 U61 (O[71], I_R[71], S);
  BWCPP_72 U62 (O[72], I_R[72], S);
  BWCPP_73 U63 (O[73], I_R[73], S);
  BWCNP_74 U64 (O[74], I_T, S);
endmodule

module TUBWCON_76_12 (O, I_T, I_R, S);
  output [76:12] O;
  input [75:12] I_R;
  input I_T;
  input S;
  BWCPP_12 U0 (O[12], I_R[12], S);
  BWCPP_13 U1 (O[13], I_R[13], S);
  BWCPP_14 U2 (O[14], I_R[14], S);
  BWCPP_15 U3 (O[15], I_R[15], S);
  BWCPP_16 U4 (O[16], I_R[16], S);
  BWCPP_17 U5 (O[17], I_R[17], S);
  BWCPP_18 U6 (O[18], I_R[18], S);
  BWCPP_19 U7 (O[19], I_R[19], S);
  BWCPP_20 U8 (O[20], I_R[20], S);
  BWCPP_21 U9 (O[21], I_R[21], S);
  BWCPP_22 U10 (O[22], I_R[22], S);
  BWCPP_23 U11 (O[23], I_R[23], S);
  BWCPP_24 U12 (O[24], I_R[24], S);
  BWCPP_25 U13 (O[25], I_R[25], S);
  BWCPP_26 U14 (O[26], I_R[26], S);
  BWCPP_27 U15 (O[27], I_R[27], S);
  BWCPP_28 U16 (O[28], I_R[28], S);
  BWCPP_29 U17 (O[29], I_R[29], S);
  BWCPP_30 U18 (O[30], I_R[30], S);
  BWCPP_31 U19 (O[31], I_R[31], S);
  BWCPP_32 U20 (O[32], I_R[32], S);
  BWCPP_33 U21 (O[33], I_R[33], S);
  BWCPP_34 U22 (O[34], I_R[34], S);
  BWCPP_35 U23 (O[35], I_R[35], S);
  BWCPP_36 U24 (O[36], I_R[36], S);
  BWCPP_37 U25 (O[37], I_R[37], S);
  BWCPP_38 U26 (O[38], I_R[38], S);
  BWCPP_39 U27 (O[39], I_R[39], S);
  BWCPP_40 U28 (O[40], I_R[40], S);
  BWCPP_41 U29 (O[41], I_R[41], S);
  BWCPP_42 U30 (O[42], I_R[42], S);
  BWCPP_43 U31 (O[43], I_R[43], S);
  BWCPP_44 U32 (O[44], I_R[44], S);
  BWCPP_45 U33 (O[45], I_R[45], S);
  BWCPP_46 U34 (O[46], I_R[46], S);
  BWCPP_47 U35 (O[47], I_R[47], S);
  BWCPP_48 U36 (O[48], I_R[48], S);
  BWCPP_49 U37 (O[49], I_R[49], S);
  BWCPP_50 U38 (O[50], I_R[50], S);
  BWCPP_51 U39 (O[51], I_R[51], S);
  BWCPP_52 U40 (O[52], I_R[52], S);
  BWCPP_53 U41 (O[53], I_R[53], S);
  BWCPP_54 U42 (O[54], I_R[54], S);
  BWCPP_55 U43 (O[55], I_R[55], S);
  BWCPP_56 U44 (O[56], I_R[56], S);
  BWCPP_57 U45 (O[57], I_R[57], S);
  BWCPP_58 U46 (O[58], I_R[58], S);
  BWCPP_59 U47 (O[59], I_R[59], S);
  BWCPP_60 U48 (O[60], I_R[60], S);
  BWCPP_61 U49 (O[61], I_R[61], S);
  BWCPP_62 U50 (O[62], I_R[62], S);
  BWCPP_63 U51 (O[63], I_R[63], S);
  BWCPP_64 U52 (O[64], I_R[64], S);
  BWCPP_65 U53 (O[65], I_R[65], S);
  BWCPP_66 U54 (O[66], I_R[66], S);
  BWCPP_67 U55 (O[67], I_R[67], S);
  BWCPP_68 U56 (O[68], I_R[68], S);
  BWCPP_69 U57 (O[69], I_R[69], S);
  BWCPP_70 U58 (O[70], I_R[70], S);
  BWCPP_71 U59 (O[71], I_R[71], S);
  BWCPP_72 U60 (O[72], I_R[72], S);
  BWCPP_73 U61 (O[73], I_R[73], S);
  BWCPP_74 U62 (O[74], I_R[74], S);
  BWCPP_75 U63 (O[75], I_R[75], S);
  BWCNP_76 U64 (O[76], I_T, S);
endmodule

module TUBWCON_78_14 (O, I_T, I_R, S);
  output [78:14] O;
  input [77:14] I_R;
  input I_T;
  input S;
  BWCPP_14 U0 (O[14], I_R[14], S);
  BWCPP_15 U1 (O[15], I_R[15], S);
  BWCPP_16 U2 (O[16], I_R[16], S);
  BWCPP_17 U3 (O[17], I_R[17], S);
  BWCPP_18 U4 (O[18], I_R[18], S);
  BWCPP_19 U5 (O[19], I_R[19], S);
  BWCPP_20 U6 (O[20], I_R[20], S);
  BWCPP_21 U7 (O[21], I_R[21], S);
  BWCPP_22 U8 (O[22], I_R[22], S);
  BWCPP_23 U9 (O[23], I_R[23], S);
  BWCPP_24 U10 (O[24], I_R[24], S);
  BWCPP_25 U11 (O[25], I_R[25], S);
  BWCPP_26 U12 (O[26], I_R[26], S);
  BWCPP_27 U13 (O[27], I_R[27], S);
  BWCPP_28 U14 (O[28], I_R[28], S);
  BWCPP_29 U15 (O[29], I_R[29], S);
  BWCPP_30 U16 (O[30], I_R[30], S);
  BWCPP_31 U17 (O[31], I_R[31], S);
  BWCPP_32 U18 (O[32], I_R[32], S);
  BWCPP_33 U19 (O[33], I_R[33], S);
  BWCPP_34 U20 (O[34], I_R[34], S);
  BWCPP_35 U21 (O[35], I_R[35], S);
  BWCPP_36 U22 (O[36], I_R[36], S);
  BWCPP_37 U23 (O[37], I_R[37], S);
  BWCPP_38 U24 (O[38], I_R[38], S);
  BWCPP_39 U25 (O[39], I_R[39], S);
  BWCPP_40 U26 (O[40], I_R[40], S);
  BWCPP_41 U27 (O[41], I_R[41], S);
  BWCPP_42 U28 (O[42], I_R[42], S);
  BWCPP_43 U29 (O[43], I_R[43], S);
  BWCPP_44 U30 (O[44], I_R[44], S);
  BWCPP_45 U31 (O[45], I_R[45], S);
  BWCPP_46 U32 (O[46], I_R[46], S);
  BWCPP_47 U33 (O[47], I_R[47], S);
  BWCPP_48 U34 (O[48], I_R[48], S);
  BWCPP_49 U35 (O[49], I_R[49], S);
  BWCPP_50 U36 (O[50], I_R[50], S);
  BWCPP_51 U37 (O[51], I_R[51], S);
  BWCPP_52 U38 (O[52], I_R[52], S);
  BWCPP_53 U39 (O[53], I_R[53], S);
  BWCPP_54 U40 (O[54], I_R[54], S);
  BWCPP_55 U41 (O[55], I_R[55], S);
  BWCPP_56 U42 (O[56], I_R[56], S);
  BWCPP_57 U43 (O[57], I_R[57], S);
  BWCPP_58 U44 (O[58], I_R[58], S);
  BWCPP_59 U45 (O[59], I_R[59], S);
  BWCPP_60 U46 (O[60], I_R[60], S);
  BWCPP_61 U47 (O[61], I_R[61], S);
  BWCPP_62 U48 (O[62], I_R[62], S);
  BWCPP_63 U49 (O[63], I_R[63], S);
  BWCPP_64 U50 (O[64], I_R[64], S);
  BWCPP_65 U51 (O[65], I_R[65], S);
  BWCPP_66 U52 (O[66], I_R[66], S);
  BWCPP_67 U53 (O[67], I_R[67], S);
  BWCPP_68 U54 (O[68], I_R[68], S);
  BWCPP_69 U55 (O[69], I_R[69], S);
  BWCPP_70 U56 (O[70], I_R[70], S);
  BWCPP_71 U57 (O[71], I_R[71], S);
  BWCPP_72 U58 (O[72], I_R[72], S);
  BWCPP_73 U59 (O[73], I_R[73], S);
  BWCPP_74 U60 (O[74], I_R[74], S);
  BWCPP_75 U61 (O[75], I_R[75], S);
  BWCPP_76 U62 (O[76], I_R[76], S);
  BWCPP_77 U63 (O[77], I_R[77], S);
  BWCNP_78 U64 (O[78], I_T, S);
endmodule

module TUBWCON_80_16 (O, I_T, I_R, S);
  output [80:16] O;
  input [79:16] I_R;
  input I_T;
  input S;
  BWCPP_16 U0 (O[16], I_R[16], S);
  BWCPP_17 U1 (O[17], I_R[17], S);
  BWCPP_18 U2 (O[18], I_R[18], S);
  BWCPP_19 U3 (O[19], I_R[19], S);
  BWCPP_20 U4 (O[20], I_R[20], S);
  BWCPP_21 U5 (O[21], I_R[21], S);
  BWCPP_22 U6 (O[22], I_R[22], S);
  BWCPP_23 U7 (O[23], I_R[23], S);
  BWCPP_24 U8 (O[24], I_R[24], S);
  BWCPP_25 U9 (O[25], I_R[25], S);
  BWCPP_26 U10 (O[26], I_R[26], S);
  BWCPP_27 U11 (O[27], I_R[27], S);
  BWCPP_28 U12 (O[28], I_R[28], S);
  BWCPP_29 U13 (O[29], I_R[29], S);
  BWCPP_30 U14 (O[30], I_R[30], S);
  BWCPP_31 U15 (O[31], I_R[31], S);
  BWCPP_32 U16 (O[32], I_R[32], S);
  BWCPP_33 U17 (O[33], I_R[33], S);
  BWCPP_34 U18 (O[34], I_R[34], S);
  BWCPP_35 U19 (O[35], I_R[35], S);
  BWCPP_36 U20 (O[36], I_R[36], S);
  BWCPP_37 U21 (O[37], I_R[37], S);
  BWCPP_38 U22 (O[38], I_R[38], S);
  BWCPP_39 U23 (O[39], I_R[39], S);
  BWCPP_40 U24 (O[40], I_R[40], S);
  BWCPP_41 U25 (O[41], I_R[41], S);
  BWCPP_42 U26 (O[42], I_R[42], S);
  BWCPP_43 U27 (O[43], I_R[43], S);
  BWCPP_44 U28 (O[44], I_R[44], S);
  BWCPP_45 U29 (O[45], I_R[45], S);
  BWCPP_46 U30 (O[46], I_R[46], S);
  BWCPP_47 U31 (O[47], I_R[47], S);
  BWCPP_48 U32 (O[48], I_R[48], S);
  BWCPP_49 U33 (O[49], I_R[49], S);
  BWCPP_50 U34 (O[50], I_R[50], S);
  BWCPP_51 U35 (O[51], I_R[51], S);
  BWCPP_52 U36 (O[52], I_R[52], S);
  BWCPP_53 U37 (O[53], I_R[53], S);
  BWCPP_54 U38 (O[54], I_R[54], S);
  BWCPP_55 U39 (O[55], I_R[55], S);
  BWCPP_56 U40 (O[56], I_R[56], S);
  BWCPP_57 U41 (O[57], I_R[57], S);
  BWCPP_58 U42 (O[58], I_R[58], S);
  BWCPP_59 U43 (O[59], I_R[59], S);
  BWCPP_60 U44 (O[60], I_R[60], S);
  BWCPP_61 U45 (O[61], I_R[61], S);
  BWCPP_62 U46 (O[62], I_R[62], S);
  BWCPP_63 U47 (O[63], I_R[63], S);
  BWCPP_64 U48 (O[64], I_R[64], S);
  BWCPP_65 U49 (O[65], I_R[65], S);
  BWCPP_66 U50 (O[66], I_R[66], S);
  BWCPP_67 U51 (O[67], I_R[67], S);
  BWCPP_68 U52 (O[68], I_R[68], S);
  BWCPP_69 U53 (O[69], I_R[69], S);
  BWCPP_70 U54 (O[70], I_R[70], S);
  BWCPP_71 U55 (O[71], I_R[71], S);
  BWCPP_72 U56 (O[72], I_R[72], S);
  BWCPP_73 U57 (O[73], I_R[73], S);
  BWCPP_74 U58 (O[74], I_R[74], S);
  BWCPP_75 U59 (O[75], I_R[75], S);
  BWCPP_76 U60 (O[76], I_R[76], S);
  BWCPP_77 U61 (O[77], I_R[77], S);
  BWCPP_78 U62 (O[78], I_R[78], S);
  BWCPP_79 U63 (O[79], I_R[79], S);
  BWCNP_80 U64 (O[80], I_T, S);
endmodule

module TUBWCON_82_18 (O, I_T, I_R, S);
  output [82:18] O;
  input [81:18] I_R;
  input I_T;
  input S;
  BWCPP_18 U0 (O[18], I_R[18], S);
  BWCPP_19 U1 (O[19], I_R[19], S);
  BWCPP_20 U2 (O[20], I_R[20], S);
  BWCPP_21 U3 (O[21], I_R[21], S);
  BWCPP_22 U4 (O[22], I_R[22], S);
  BWCPP_23 U5 (O[23], I_R[23], S);
  BWCPP_24 U6 (O[24], I_R[24], S);
  BWCPP_25 U7 (O[25], I_R[25], S);
  BWCPP_26 U8 (O[26], I_R[26], S);
  BWCPP_27 U9 (O[27], I_R[27], S);
  BWCPP_28 U10 (O[28], I_R[28], S);
  BWCPP_29 U11 (O[29], I_R[29], S);
  BWCPP_30 U12 (O[30], I_R[30], S);
  BWCPP_31 U13 (O[31], I_R[31], S);
  BWCPP_32 U14 (O[32], I_R[32], S);
  BWCPP_33 U15 (O[33], I_R[33], S);
  BWCPP_34 U16 (O[34], I_R[34], S);
  BWCPP_35 U17 (O[35], I_R[35], S);
  BWCPP_36 U18 (O[36], I_R[36], S);
  BWCPP_37 U19 (O[37], I_R[37], S);
  BWCPP_38 U20 (O[38], I_R[38], S);
  BWCPP_39 U21 (O[39], I_R[39], S);
  BWCPP_40 U22 (O[40], I_R[40], S);
  BWCPP_41 U23 (O[41], I_R[41], S);
  BWCPP_42 U24 (O[42], I_R[42], S);
  BWCPP_43 U25 (O[43], I_R[43], S);
  BWCPP_44 U26 (O[44], I_R[44], S);
  BWCPP_45 U27 (O[45], I_R[45], S);
  BWCPP_46 U28 (O[46], I_R[46], S);
  BWCPP_47 U29 (O[47], I_R[47], S);
  BWCPP_48 U30 (O[48], I_R[48], S);
  BWCPP_49 U31 (O[49], I_R[49], S);
  BWCPP_50 U32 (O[50], I_R[50], S);
  BWCPP_51 U33 (O[51], I_R[51], S);
  BWCPP_52 U34 (O[52], I_R[52], S);
  BWCPP_53 U35 (O[53], I_R[53], S);
  BWCPP_54 U36 (O[54], I_R[54], S);
  BWCPP_55 U37 (O[55], I_R[55], S);
  BWCPP_56 U38 (O[56], I_R[56], S);
  BWCPP_57 U39 (O[57], I_R[57], S);
  BWCPP_58 U40 (O[58], I_R[58], S);
  BWCPP_59 U41 (O[59], I_R[59], S);
  BWCPP_60 U42 (O[60], I_R[60], S);
  BWCPP_61 U43 (O[61], I_R[61], S);
  BWCPP_62 U44 (O[62], I_R[62], S);
  BWCPP_63 U45 (O[63], I_R[63], S);
  BWCPP_64 U46 (O[64], I_R[64], S);
  BWCPP_65 U47 (O[65], I_R[65], S);
  BWCPP_66 U48 (O[66], I_R[66], S);
  BWCPP_67 U49 (O[67], I_R[67], S);
  BWCPP_68 U50 (O[68], I_R[68], S);
  BWCPP_69 U51 (O[69], I_R[69], S);
  BWCPP_70 U52 (O[70], I_R[70], S);
  BWCPP_71 U53 (O[71], I_R[71], S);
  BWCPP_72 U54 (O[72], I_R[72], S);
  BWCPP_73 U55 (O[73], I_R[73], S);
  BWCPP_74 U56 (O[74], I_R[74], S);
  BWCPP_75 U57 (O[75], I_R[75], S);
  BWCPP_76 U58 (O[76], I_R[76], S);
  BWCPP_77 U59 (O[77], I_R[77], S);
  BWCPP_78 U60 (O[78], I_R[78], S);
  BWCPP_79 U61 (O[79], I_R[79], S);
  BWCPP_80 U62 (O[80], I_R[80], S);
  BWCPP_81 U63 (O[81], I_R[81], S);
  BWCNP_82 U64 (O[82], I_T, S);
endmodule

module TUBWCON_84_20 (O, I_T, I_R, S);
  output [84:20] O;
  input [83:20] I_R;
  input I_T;
  input S;
  BWCPP_20 U0 (O[20], I_R[20], S);
  BWCPP_21 U1 (O[21], I_R[21], S);
  BWCPP_22 U2 (O[22], I_R[22], S);
  BWCPP_23 U3 (O[23], I_R[23], S);
  BWCPP_24 U4 (O[24], I_R[24], S);
  BWCPP_25 U5 (O[25], I_R[25], S);
  BWCPP_26 U6 (O[26], I_R[26], S);
  BWCPP_27 U7 (O[27], I_R[27], S);
  BWCPP_28 U8 (O[28], I_R[28], S);
  BWCPP_29 U9 (O[29], I_R[29], S);
  BWCPP_30 U10 (O[30], I_R[30], S);
  BWCPP_31 U11 (O[31], I_R[31], S);
  BWCPP_32 U12 (O[32], I_R[32], S);
  BWCPP_33 U13 (O[33], I_R[33], S);
  BWCPP_34 U14 (O[34], I_R[34], S);
  BWCPP_35 U15 (O[35], I_R[35], S);
  BWCPP_36 U16 (O[36], I_R[36], S);
  BWCPP_37 U17 (O[37], I_R[37], S);
  BWCPP_38 U18 (O[38], I_R[38], S);
  BWCPP_39 U19 (O[39], I_R[39], S);
  BWCPP_40 U20 (O[40], I_R[40], S);
  BWCPP_41 U21 (O[41], I_R[41], S);
  BWCPP_42 U22 (O[42], I_R[42], S);
  BWCPP_43 U23 (O[43], I_R[43], S);
  BWCPP_44 U24 (O[44], I_R[44], S);
  BWCPP_45 U25 (O[45], I_R[45], S);
  BWCPP_46 U26 (O[46], I_R[46], S);
  BWCPP_47 U27 (O[47], I_R[47], S);
  BWCPP_48 U28 (O[48], I_R[48], S);
  BWCPP_49 U29 (O[49], I_R[49], S);
  BWCPP_50 U30 (O[50], I_R[50], S);
  BWCPP_51 U31 (O[51], I_R[51], S);
  BWCPP_52 U32 (O[52], I_R[52], S);
  BWCPP_53 U33 (O[53], I_R[53], S);
  BWCPP_54 U34 (O[54], I_R[54], S);
  BWCPP_55 U35 (O[55], I_R[55], S);
  BWCPP_56 U36 (O[56], I_R[56], S);
  BWCPP_57 U37 (O[57], I_R[57], S);
  BWCPP_58 U38 (O[58], I_R[58], S);
  BWCPP_59 U39 (O[59], I_R[59], S);
  BWCPP_60 U40 (O[60], I_R[60], S);
  BWCPP_61 U41 (O[61], I_R[61], S);
  BWCPP_62 U42 (O[62], I_R[62], S);
  BWCPP_63 U43 (O[63], I_R[63], S);
  BWCPP_64 U44 (O[64], I_R[64], S);
  BWCPP_65 U45 (O[65], I_R[65], S);
  BWCPP_66 U46 (O[66], I_R[66], S);
  BWCPP_67 U47 (O[67], I_R[67], S);
  BWCPP_68 U48 (O[68], I_R[68], S);
  BWCPP_69 U49 (O[69], I_R[69], S);
  BWCPP_70 U50 (O[70], I_R[70], S);
  BWCPP_71 U51 (O[71], I_R[71], S);
  BWCPP_72 U52 (O[72], I_R[72], S);
  BWCPP_73 U53 (O[73], I_R[73], S);
  BWCPP_74 U54 (O[74], I_R[74], S);
  BWCPP_75 U55 (O[75], I_R[75], S);
  BWCPP_76 U56 (O[76], I_R[76], S);
  BWCPP_77 U57 (O[77], I_R[77], S);
  BWCPP_78 U58 (O[78], I_R[78], S);
  BWCPP_79 U59 (O[79], I_R[79], S);
  BWCPP_80 U60 (O[80], I_R[80], S);
  BWCPP_81 U61 (O[81], I_R[81], S);
  BWCPP_82 U62 (O[82], I_R[82], S);
  BWCPP_83 U63 (O[83], I_R[83], S);
  BWCNP_84 U64 (O[84], I_T, S);
endmodule

module TUBWCON_86_22 (O, I_T, I_R, S);
  output [86:22] O;
  input [85:22] I_R;
  input I_T;
  input S;
  BWCPP_22 U0 (O[22], I_R[22], S);
  BWCPP_23 U1 (O[23], I_R[23], S);
  BWCPP_24 U2 (O[24], I_R[24], S);
  BWCPP_25 U3 (O[25], I_R[25], S);
  BWCPP_26 U4 (O[26], I_R[26], S);
  BWCPP_27 U5 (O[27], I_R[27], S);
  BWCPP_28 U6 (O[28], I_R[28], S);
  BWCPP_29 U7 (O[29], I_R[29], S);
  BWCPP_30 U8 (O[30], I_R[30], S);
  BWCPP_31 U9 (O[31], I_R[31], S);
  BWCPP_32 U10 (O[32], I_R[32], S);
  BWCPP_33 U11 (O[33], I_R[33], S);
  BWCPP_34 U12 (O[34], I_R[34], S);
  BWCPP_35 U13 (O[35], I_R[35], S);
  BWCPP_36 U14 (O[36], I_R[36], S);
  BWCPP_37 U15 (O[37], I_R[37], S);
  BWCPP_38 U16 (O[38], I_R[38], S);
  BWCPP_39 U17 (O[39], I_R[39], S);
  BWCPP_40 U18 (O[40], I_R[40], S);
  BWCPP_41 U19 (O[41], I_R[41], S);
  BWCPP_42 U20 (O[42], I_R[42], S);
  BWCPP_43 U21 (O[43], I_R[43], S);
  BWCPP_44 U22 (O[44], I_R[44], S);
  BWCPP_45 U23 (O[45], I_R[45], S);
  BWCPP_46 U24 (O[46], I_R[46], S);
  BWCPP_47 U25 (O[47], I_R[47], S);
  BWCPP_48 U26 (O[48], I_R[48], S);
  BWCPP_49 U27 (O[49], I_R[49], S);
  BWCPP_50 U28 (O[50], I_R[50], S);
  BWCPP_51 U29 (O[51], I_R[51], S);
  BWCPP_52 U30 (O[52], I_R[52], S);
  BWCPP_53 U31 (O[53], I_R[53], S);
  BWCPP_54 U32 (O[54], I_R[54], S);
  BWCPP_55 U33 (O[55], I_R[55], S);
  BWCPP_56 U34 (O[56], I_R[56], S);
  BWCPP_57 U35 (O[57], I_R[57], S);
  BWCPP_58 U36 (O[58], I_R[58], S);
  BWCPP_59 U37 (O[59], I_R[59], S);
  BWCPP_60 U38 (O[60], I_R[60], S);
  BWCPP_61 U39 (O[61], I_R[61], S);
  BWCPP_62 U40 (O[62], I_R[62], S);
  BWCPP_63 U41 (O[63], I_R[63], S);
  BWCPP_64 U42 (O[64], I_R[64], S);
  BWCPP_65 U43 (O[65], I_R[65], S);
  BWCPP_66 U44 (O[66], I_R[66], S);
  BWCPP_67 U45 (O[67], I_R[67], S);
  BWCPP_68 U46 (O[68], I_R[68], S);
  BWCPP_69 U47 (O[69], I_R[69], S);
  BWCPP_70 U48 (O[70], I_R[70], S);
  BWCPP_71 U49 (O[71], I_R[71], S);
  BWCPP_72 U50 (O[72], I_R[72], S);
  BWCPP_73 U51 (O[73], I_R[73], S);
  BWCPP_74 U52 (O[74], I_R[74], S);
  BWCPP_75 U53 (O[75], I_R[75], S);
  BWCPP_76 U54 (O[76], I_R[76], S);
  BWCPP_77 U55 (O[77], I_R[77], S);
  BWCPP_78 U56 (O[78], I_R[78], S);
  BWCPP_79 U57 (O[79], I_R[79], S);
  BWCPP_80 U58 (O[80], I_R[80], S);
  BWCPP_81 U59 (O[81], I_R[81], S);
  BWCPP_82 U60 (O[82], I_R[82], S);
  BWCPP_83 U61 (O[83], I_R[83], S);
  BWCPP_84 U62 (O[84], I_R[84], S);
  BWCPP_85 U63 (O[85], I_R[85], S);
  BWCNP_86 U64 (O[86], I_T, S);
endmodule

module TUBWCON_88_24 (O, I_T, I_R, S);
  output [88:24] O;
  input [87:24] I_R;
  input I_T;
  input S;
  BWCPP_24 U0 (O[24], I_R[24], S);
  BWCPP_25 U1 (O[25], I_R[25], S);
  BWCPP_26 U2 (O[26], I_R[26], S);
  BWCPP_27 U3 (O[27], I_R[27], S);
  BWCPP_28 U4 (O[28], I_R[28], S);
  BWCPP_29 U5 (O[29], I_R[29], S);
  BWCPP_30 U6 (O[30], I_R[30], S);
  BWCPP_31 U7 (O[31], I_R[31], S);
  BWCPP_32 U8 (O[32], I_R[32], S);
  BWCPP_33 U9 (O[33], I_R[33], S);
  BWCPP_34 U10 (O[34], I_R[34], S);
  BWCPP_35 U11 (O[35], I_R[35], S);
  BWCPP_36 U12 (O[36], I_R[36], S);
  BWCPP_37 U13 (O[37], I_R[37], S);
  BWCPP_38 U14 (O[38], I_R[38], S);
  BWCPP_39 U15 (O[39], I_R[39], S);
  BWCPP_40 U16 (O[40], I_R[40], S);
  BWCPP_41 U17 (O[41], I_R[41], S);
  BWCPP_42 U18 (O[42], I_R[42], S);
  BWCPP_43 U19 (O[43], I_R[43], S);
  BWCPP_44 U20 (O[44], I_R[44], S);
  BWCPP_45 U21 (O[45], I_R[45], S);
  BWCPP_46 U22 (O[46], I_R[46], S);
  BWCPP_47 U23 (O[47], I_R[47], S);
  BWCPP_48 U24 (O[48], I_R[48], S);
  BWCPP_49 U25 (O[49], I_R[49], S);
  BWCPP_50 U26 (O[50], I_R[50], S);
  BWCPP_51 U27 (O[51], I_R[51], S);
  BWCPP_52 U28 (O[52], I_R[52], S);
  BWCPP_53 U29 (O[53], I_R[53], S);
  BWCPP_54 U30 (O[54], I_R[54], S);
  BWCPP_55 U31 (O[55], I_R[55], S);
  BWCPP_56 U32 (O[56], I_R[56], S);
  BWCPP_57 U33 (O[57], I_R[57], S);
  BWCPP_58 U34 (O[58], I_R[58], S);
  BWCPP_59 U35 (O[59], I_R[59], S);
  BWCPP_60 U36 (O[60], I_R[60], S);
  BWCPP_61 U37 (O[61], I_R[61], S);
  BWCPP_62 U38 (O[62], I_R[62], S);
  BWCPP_63 U39 (O[63], I_R[63], S);
  BWCPP_64 U40 (O[64], I_R[64], S);
  BWCPP_65 U41 (O[65], I_R[65], S);
  BWCPP_66 U42 (O[66], I_R[66], S);
  BWCPP_67 U43 (O[67], I_R[67], S);
  BWCPP_68 U44 (O[68], I_R[68], S);
  BWCPP_69 U45 (O[69], I_R[69], S);
  BWCPP_70 U46 (O[70], I_R[70], S);
  BWCPP_71 U47 (O[71], I_R[71], S);
  BWCPP_72 U48 (O[72], I_R[72], S);
  BWCPP_73 U49 (O[73], I_R[73], S);
  BWCPP_74 U50 (O[74], I_R[74], S);
  BWCPP_75 U51 (O[75], I_R[75], S);
  BWCPP_76 U52 (O[76], I_R[76], S);
  BWCPP_77 U53 (O[77], I_R[77], S);
  BWCPP_78 U54 (O[78], I_R[78], S);
  BWCPP_79 U55 (O[79], I_R[79], S);
  BWCPP_80 U56 (O[80], I_R[80], S);
  BWCPP_81 U57 (O[81], I_R[81], S);
  BWCPP_82 U58 (O[82], I_R[82], S);
  BWCPP_83 U59 (O[83], I_R[83], S);
  BWCPP_84 U60 (O[84], I_R[84], S);
  BWCPP_85 U61 (O[85], I_R[85], S);
  BWCPP_86 U62 (O[86], I_R[86], S);
  BWCPP_87 U63 (O[87], I_R[87], S);
  BWCNP_88 U64 (O[88], I_T, S);
endmodule

module TUBWCON_90_26 (O, I_T, I_R, S);
  output [90:26] O;
  input [89:26] I_R;
  input I_T;
  input S;
  BWCPP_26 U0 (O[26], I_R[26], S);
  BWCPP_27 U1 (O[27], I_R[27], S);
  BWCPP_28 U2 (O[28], I_R[28], S);
  BWCPP_29 U3 (O[29], I_R[29], S);
  BWCPP_30 U4 (O[30], I_R[30], S);
  BWCPP_31 U5 (O[31], I_R[31], S);
  BWCPP_32 U6 (O[32], I_R[32], S);
  BWCPP_33 U7 (O[33], I_R[33], S);
  BWCPP_34 U8 (O[34], I_R[34], S);
  BWCPP_35 U9 (O[35], I_R[35], S);
  BWCPP_36 U10 (O[36], I_R[36], S);
  BWCPP_37 U11 (O[37], I_R[37], S);
  BWCPP_38 U12 (O[38], I_R[38], S);
  BWCPP_39 U13 (O[39], I_R[39], S);
  BWCPP_40 U14 (O[40], I_R[40], S);
  BWCPP_41 U15 (O[41], I_R[41], S);
  BWCPP_42 U16 (O[42], I_R[42], S);
  BWCPP_43 U17 (O[43], I_R[43], S);
  BWCPP_44 U18 (O[44], I_R[44], S);
  BWCPP_45 U19 (O[45], I_R[45], S);
  BWCPP_46 U20 (O[46], I_R[46], S);
  BWCPP_47 U21 (O[47], I_R[47], S);
  BWCPP_48 U22 (O[48], I_R[48], S);
  BWCPP_49 U23 (O[49], I_R[49], S);
  BWCPP_50 U24 (O[50], I_R[50], S);
  BWCPP_51 U25 (O[51], I_R[51], S);
  BWCPP_52 U26 (O[52], I_R[52], S);
  BWCPP_53 U27 (O[53], I_R[53], S);
  BWCPP_54 U28 (O[54], I_R[54], S);
  BWCPP_55 U29 (O[55], I_R[55], S);
  BWCPP_56 U30 (O[56], I_R[56], S);
  BWCPP_57 U31 (O[57], I_R[57], S);
  BWCPP_58 U32 (O[58], I_R[58], S);
  BWCPP_59 U33 (O[59], I_R[59], S);
  BWCPP_60 U34 (O[60], I_R[60], S);
  BWCPP_61 U35 (O[61], I_R[61], S);
  BWCPP_62 U36 (O[62], I_R[62], S);
  BWCPP_63 U37 (O[63], I_R[63], S);
  BWCPP_64 U38 (O[64], I_R[64], S);
  BWCPP_65 U39 (O[65], I_R[65], S);
  BWCPP_66 U40 (O[66], I_R[66], S);
  BWCPP_67 U41 (O[67], I_R[67], S);
  BWCPP_68 U42 (O[68], I_R[68], S);
  BWCPP_69 U43 (O[69], I_R[69], S);
  BWCPP_70 U44 (O[70], I_R[70], S);
  BWCPP_71 U45 (O[71], I_R[71], S);
  BWCPP_72 U46 (O[72], I_R[72], S);
  BWCPP_73 U47 (O[73], I_R[73], S);
  BWCPP_74 U48 (O[74], I_R[74], S);
  BWCPP_75 U49 (O[75], I_R[75], S);
  BWCPP_76 U50 (O[76], I_R[76], S);
  BWCPP_77 U51 (O[77], I_R[77], S);
  BWCPP_78 U52 (O[78], I_R[78], S);
  BWCPP_79 U53 (O[79], I_R[79], S);
  BWCPP_80 U54 (O[80], I_R[80], S);
  BWCPP_81 U55 (O[81], I_R[81], S);
  BWCPP_82 U56 (O[82], I_R[82], S);
  BWCPP_83 U57 (O[83], I_R[83], S);
  BWCPP_84 U58 (O[84], I_R[84], S);
  BWCPP_85 U59 (O[85], I_R[85], S);
  BWCPP_86 U60 (O[86], I_R[86], S);
  BWCPP_87 U61 (O[87], I_R[87], S);
  BWCPP_88 U62 (O[88], I_R[88], S);
  BWCPP_89 U63 (O[89], I_R[89], S);
  BWCNP_90 U64 (O[90], I_T, S);
endmodule

module TUBWCON_92_28 (O, I_T, I_R, S);
  output [92:28] O;
  input [91:28] I_R;
  input I_T;
  input S;
  BWCPP_28 U0 (O[28], I_R[28], S);
  BWCPP_29 U1 (O[29], I_R[29], S);
  BWCPP_30 U2 (O[30], I_R[30], S);
  BWCPP_31 U3 (O[31], I_R[31], S);
  BWCPP_32 U4 (O[32], I_R[32], S);
  BWCPP_33 U5 (O[33], I_R[33], S);
  BWCPP_34 U6 (O[34], I_R[34], S);
  BWCPP_35 U7 (O[35], I_R[35], S);
  BWCPP_36 U8 (O[36], I_R[36], S);
  BWCPP_37 U9 (O[37], I_R[37], S);
  BWCPP_38 U10 (O[38], I_R[38], S);
  BWCPP_39 U11 (O[39], I_R[39], S);
  BWCPP_40 U12 (O[40], I_R[40], S);
  BWCPP_41 U13 (O[41], I_R[41], S);
  BWCPP_42 U14 (O[42], I_R[42], S);
  BWCPP_43 U15 (O[43], I_R[43], S);
  BWCPP_44 U16 (O[44], I_R[44], S);
  BWCPP_45 U17 (O[45], I_R[45], S);
  BWCPP_46 U18 (O[46], I_R[46], S);
  BWCPP_47 U19 (O[47], I_R[47], S);
  BWCPP_48 U20 (O[48], I_R[48], S);
  BWCPP_49 U21 (O[49], I_R[49], S);
  BWCPP_50 U22 (O[50], I_R[50], S);
  BWCPP_51 U23 (O[51], I_R[51], S);
  BWCPP_52 U24 (O[52], I_R[52], S);
  BWCPP_53 U25 (O[53], I_R[53], S);
  BWCPP_54 U26 (O[54], I_R[54], S);
  BWCPP_55 U27 (O[55], I_R[55], S);
  BWCPP_56 U28 (O[56], I_R[56], S);
  BWCPP_57 U29 (O[57], I_R[57], S);
  BWCPP_58 U30 (O[58], I_R[58], S);
  BWCPP_59 U31 (O[59], I_R[59], S);
  BWCPP_60 U32 (O[60], I_R[60], S);
  BWCPP_61 U33 (O[61], I_R[61], S);
  BWCPP_62 U34 (O[62], I_R[62], S);
  BWCPP_63 U35 (O[63], I_R[63], S);
  BWCPP_64 U36 (O[64], I_R[64], S);
  BWCPP_65 U37 (O[65], I_R[65], S);
  BWCPP_66 U38 (O[66], I_R[66], S);
  BWCPP_67 U39 (O[67], I_R[67], S);
  BWCPP_68 U40 (O[68], I_R[68], S);
  BWCPP_69 U41 (O[69], I_R[69], S);
  BWCPP_70 U42 (O[70], I_R[70], S);
  BWCPP_71 U43 (O[71], I_R[71], S);
  BWCPP_72 U44 (O[72], I_R[72], S);
  BWCPP_73 U45 (O[73], I_R[73], S);
  BWCPP_74 U46 (O[74], I_R[74], S);
  BWCPP_75 U47 (O[75], I_R[75], S);
  BWCPP_76 U48 (O[76], I_R[76], S);
  BWCPP_77 U49 (O[77], I_R[77], S);
  BWCPP_78 U50 (O[78], I_R[78], S);
  BWCPP_79 U51 (O[79], I_R[79], S);
  BWCPP_80 U52 (O[80], I_R[80], S);
  BWCPP_81 U53 (O[81], I_R[81], S);
  BWCPP_82 U54 (O[82], I_R[82], S);
  BWCPP_83 U55 (O[83], I_R[83], S);
  BWCPP_84 U56 (O[84], I_R[84], S);
  BWCPP_85 U57 (O[85], I_R[85], S);
  BWCPP_86 U58 (O[86], I_R[86], S);
  BWCPP_87 U59 (O[87], I_R[87], S);
  BWCPP_88 U60 (O[88], I_R[88], S);
  BWCPP_89 U61 (O[89], I_R[89], S);
  BWCPP_90 U62 (O[90], I_R[90], S);
  BWCPP_91 U63 (O[91], I_R[91], S);
  BWCNP_92 U64 (O[92], I_T, S);
endmodule

module TUBWCON_94_30 (O, I_T, I_R, S);
  output [94:30] O;
  input [93:30] I_R;
  input I_T;
  input S;
  BWCPP_30 U0 (O[30], I_R[30], S);
  BWCPP_31 U1 (O[31], I_R[31], S);
  BWCPP_32 U2 (O[32], I_R[32], S);
  BWCPP_33 U3 (O[33], I_R[33], S);
  BWCPP_34 U4 (O[34], I_R[34], S);
  BWCPP_35 U5 (O[35], I_R[35], S);
  BWCPP_36 U6 (O[36], I_R[36], S);
  BWCPP_37 U7 (O[37], I_R[37], S);
  BWCPP_38 U8 (O[38], I_R[38], S);
  BWCPP_39 U9 (O[39], I_R[39], S);
  BWCPP_40 U10 (O[40], I_R[40], S);
  BWCPP_41 U11 (O[41], I_R[41], S);
  BWCPP_42 U12 (O[42], I_R[42], S);
  BWCPP_43 U13 (O[43], I_R[43], S);
  BWCPP_44 U14 (O[44], I_R[44], S);
  BWCPP_45 U15 (O[45], I_R[45], S);
  BWCPP_46 U16 (O[46], I_R[46], S);
  BWCPP_47 U17 (O[47], I_R[47], S);
  BWCPP_48 U18 (O[48], I_R[48], S);
  BWCPP_49 U19 (O[49], I_R[49], S);
  BWCPP_50 U20 (O[50], I_R[50], S);
  BWCPP_51 U21 (O[51], I_R[51], S);
  BWCPP_52 U22 (O[52], I_R[52], S);
  BWCPP_53 U23 (O[53], I_R[53], S);
  BWCPP_54 U24 (O[54], I_R[54], S);
  BWCPP_55 U25 (O[55], I_R[55], S);
  BWCPP_56 U26 (O[56], I_R[56], S);
  BWCPP_57 U27 (O[57], I_R[57], S);
  BWCPP_58 U28 (O[58], I_R[58], S);
  BWCPP_59 U29 (O[59], I_R[59], S);
  BWCPP_60 U30 (O[60], I_R[60], S);
  BWCPP_61 U31 (O[61], I_R[61], S);
  BWCPP_62 U32 (O[62], I_R[62], S);
  BWCPP_63 U33 (O[63], I_R[63], S);
  BWCPP_64 U34 (O[64], I_R[64], S);
  BWCPP_65 U35 (O[65], I_R[65], S);
  BWCPP_66 U36 (O[66], I_R[66], S);
  BWCPP_67 U37 (O[67], I_R[67], S);
  BWCPP_68 U38 (O[68], I_R[68], S);
  BWCPP_69 U39 (O[69], I_R[69], S);
  BWCPP_70 U40 (O[70], I_R[70], S);
  BWCPP_71 U41 (O[71], I_R[71], S);
  BWCPP_72 U42 (O[72], I_R[72], S);
  BWCPP_73 U43 (O[73], I_R[73], S);
  BWCPP_74 U44 (O[74], I_R[74], S);
  BWCPP_75 U45 (O[75], I_R[75], S);
  BWCPP_76 U46 (O[76], I_R[76], S);
  BWCPP_77 U47 (O[77], I_R[77], S);
  BWCPP_78 U48 (O[78], I_R[78], S);
  BWCPP_79 U49 (O[79], I_R[79], S);
  BWCPP_80 U50 (O[80], I_R[80], S);
  BWCPP_81 U51 (O[81], I_R[81], S);
  BWCPP_82 U52 (O[82], I_R[82], S);
  BWCPP_83 U53 (O[83], I_R[83], S);
  BWCPP_84 U54 (O[84], I_R[84], S);
  BWCPP_85 U55 (O[85], I_R[85], S);
  BWCPP_86 U56 (O[86], I_R[86], S);
  BWCPP_87 U57 (O[87], I_R[87], S);
  BWCPP_88 U58 (O[88], I_R[88], S);
  BWCPP_89 U59 (O[89], I_R[89], S);
  BWCPP_90 U60 (O[90], I_R[90], S);
  BWCPP_91 U61 (O[91], I_R[91], S);
  BWCPP_92 U62 (O[92], I_R[92], S);
  BWCPP_93 U63 (O[93], I_R[93], S);
  BWCNP_94 U64 (O[94], I_T, S);
endmodule

module TUBWCON_96_32 (O, I_T, I_R, S);
  output [96:32] O;
  input [95:32] I_R;
  input I_T;
  input S;
  BWCPP_32 U0 (O[32], I_R[32], S);
  BWCPP_33 U1 (O[33], I_R[33], S);
  BWCPP_34 U2 (O[34], I_R[34], S);
  BWCPP_35 U3 (O[35], I_R[35], S);
  BWCPP_36 U4 (O[36], I_R[36], S);
  BWCPP_37 U5 (O[37], I_R[37], S);
  BWCPP_38 U6 (O[38], I_R[38], S);
  BWCPP_39 U7 (O[39], I_R[39], S);
  BWCPP_40 U8 (O[40], I_R[40], S);
  BWCPP_41 U9 (O[41], I_R[41], S);
  BWCPP_42 U10 (O[42], I_R[42], S);
  BWCPP_43 U11 (O[43], I_R[43], S);
  BWCPP_44 U12 (O[44], I_R[44], S);
  BWCPP_45 U13 (O[45], I_R[45], S);
  BWCPP_46 U14 (O[46], I_R[46], S);
  BWCPP_47 U15 (O[47], I_R[47], S);
  BWCPP_48 U16 (O[48], I_R[48], S);
  BWCPP_49 U17 (O[49], I_R[49], S);
  BWCPP_50 U18 (O[50], I_R[50], S);
  BWCPP_51 U19 (O[51], I_R[51], S);
  BWCPP_52 U20 (O[52], I_R[52], S);
  BWCPP_53 U21 (O[53], I_R[53], S);
  BWCPP_54 U22 (O[54], I_R[54], S);
  BWCPP_55 U23 (O[55], I_R[55], S);
  BWCPP_56 U24 (O[56], I_R[56], S);
  BWCPP_57 U25 (O[57], I_R[57], S);
  BWCPP_58 U26 (O[58], I_R[58], S);
  BWCPP_59 U27 (O[59], I_R[59], S);
  BWCPP_60 U28 (O[60], I_R[60], S);
  BWCPP_61 U29 (O[61], I_R[61], S);
  BWCPP_62 U30 (O[62], I_R[62], S);
  BWCPP_63 U31 (O[63], I_R[63], S);
  BWCPP_64 U32 (O[64], I_R[64], S);
  BWCPP_65 U33 (O[65], I_R[65], S);
  BWCPP_66 U34 (O[66], I_R[66], S);
  BWCPP_67 U35 (O[67], I_R[67], S);
  BWCPP_68 U36 (O[68], I_R[68], S);
  BWCPP_69 U37 (O[69], I_R[69], S);
  BWCPP_70 U38 (O[70], I_R[70], S);
  BWCPP_71 U39 (O[71], I_R[71], S);
  BWCPP_72 U40 (O[72], I_R[72], S);
  BWCPP_73 U41 (O[73], I_R[73], S);
  BWCPP_74 U42 (O[74], I_R[74], S);
  BWCPP_75 U43 (O[75], I_R[75], S);
  BWCPP_76 U44 (O[76], I_R[76], S);
  BWCPP_77 U45 (O[77], I_R[77], S);
  BWCPP_78 U46 (O[78], I_R[78], S);
  BWCPP_79 U47 (O[79], I_R[79], S);
  BWCPP_80 U48 (O[80], I_R[80], S);
  BWCPP_81 U49 (O[81], I_R[81], S);
  BWCPP_82 U50 (O[82], I_R[82], S);
  BWCPP_83 U51 (O[83], I_R[83], S);
  BWCPP_84 U52 (O[84], I_R[84], S);
  BWCPP_85 U53 (O[85], I_R[85], S);
  BWCPP_86 U54 (O[86], I_R[86], S);
  BWCPP_87 U55 (O[87], I_R[87], S);
  BWCPP_88 U56 (O[88], I_R[88], S);
  BWCPP_89 U57 (O[89], I_R[89], S);
  BWCPP_90 U58 (O[90], I_R[90], S);
  BWCPP_91 U59 (O[91], I_R[91], S);
  BWCPP_92 U60 (O[92], I_R[92], S);
  BWCPP_93 U61 (O[93], I_R[93], S);
  BWCPP_94 U62 (O[94], I_R[94], S);
  BWCPP_95 U63 (O[95], I_R[95], S);
  BWCNP_96 U64 (O[96], I_T, S);
endmodule

module TUBWCON_98_34 (O, I_T, I_R, S);
  output [98:34] O;
  input [97:34] I_R;
  input I_T;
  input S;
  BWCPP_34 U0 (O[34], I_R[34], S);
  BWCPP_35 U1 (O[35], I_R[35], S);
  BWCPP_36 U2 (O[36], I_R[36], S);
  BWCPP_37 U3 (O[37], I_R[37], S);
  BWCPP_38 U4 (O[38], I_R[38], S);
  BWCPP_39 U5 (O[39], I_R[39], S);
  BWCPP_40 U6 (O[40], I_R[40], S);
  BWCPP_41 U7 (O[41], I_R[41], S);
  BWCPP_42 U8 (O[42], I_R[42], S);
  BWCPP_43 U9 (O[43], I_R[43], S);
  BWCPP_44 U10 (O[44], I_R[44], S);
  BWCPP_45 U11 (O[45], I_R[45], S);
  BWCPP_46 U12 (O[46], I_R[46], S);
  BWCPP_47 U13 (O[47], I_R[47], S);
  BWCPP_48 U14 (O[48], I_R[48], S);
  BWCPP_49 U15 (O[49], I_R[49], S);
  BWCPP_50 U16 (O[50], I_R[50], S);
  BWCPP_51 U17 (O[51], I_R[51], S);
  BWCPP_52 U18 (O[52], I_R[52], S);
  BWCPP_53 U19 (O[53], I_R[53], S);
  BWCPP_54 U20 (O[54], I_R[54], S);
  BWCPP_55 U21 (O[55], I_R[55], S);
  BWCPP_56 U22 (O[56], I_R[56], S);
  BWCPP_57 U23 (O[57], I_R[57], S);
  BWCPP_58 U24 (O[58], I_R[58], S);
  BWCPP_59 U25 (O[59], I_R[59], S);
  BWCPP_60 U26 (O[60], I_R[60], S);
  BWCPP_61 U27 (O[61], I_R[61], S);
  BWCPP_62 U28 (O[62], I_R[62], S);
  BWCPP_63 U29 (O[63], I_R[63], S);
  BWCPP_64 U30 (O[64], I_R[64], S);
  BWCPP_65 U31 (O[65], I_R[65], S);
  BWCPP_66 U32 (O[66], I_R[66], S);
  BWCPP_67 U33 (O[67], I_R[67], S);
  BWCPP_68 U34 (O[68], I_R[68], S);
  BWCPP_69 U35 (O[69], I_R[69], S);
  BWCPP_70 U36 (O[70], I_R[70], S);
  BWCPP_71 U37 (O[71], I_R[71], S);
  BWCPP_72 U38 (O[72], I_R[72], S);
  BWCPP_73 U39 (O[73], I_R[73], S);
  BWCPP_74 U40 (O[74], I_R[74], S);
  BWCPP_75 U41 (O[75], I_R[75], S);
  BWCPP_76 U42 (O[76], I_R[76], S);
  BWCPP_77 U43 (O[77], I_R[77], S);
  BWCPP_78 U44 (O[78], I_R[78], S);
  BWCPP_79 U45 (O[79], I_R[79], S);
  BWCPP_80 U46 (O[80], I_R[80], S);
  BWCPP_81 U47 (O[81], I_R[81], S);
  BWCPP_82 U48 (O[82], I_R[82], S);
  BWCPP_83 U49 (O[83], I_R[83], S);
  BWCPP_84 U50 (O[84], I_R[84], S);
  BWCPP_85 U51 (O[85], I_R[85], S);
  BWCPP_86 U52 (O[86], I_R[86], S);
  BWCPP_87 U53 (O[87], I_R[87], S);
  BWCPP_88 U54 (O[88], I_R[88], S);
  BWCPP_89 U55 (O[89], I_R[89], S);
  BWCPP_90 U56 (O[90], I_R[90], S);
  BWCPP_91 U57 (O[91], I_R[91], S);
  BWCPP_92 U58 (O[92], I_R[92], S);
  BWCPP_93 U59 (O[93], I_R[93], S);
  BWCPP_94 U60 (O[94], I_R[94], S);
  BWCPP_95 U61 (O[95], I_R[95], S);
  BWCPP_96 U62 (O[96], I_R[96], S);
  BWCPP_97 U63 (O[97], I_R[97], S);
  BWCNP_98 U64 (O[98], I_T, S);
endmodule

module UBCMBIN_101_101_1000 (O, IN0, IN1, IN2);
  output [101:34] O;
  input IN0;
  input [100:36] IN1;
  input IN2;
  UB1DCON_101 U0 (O[101], IN0);
  UBCON_100_36 U1 (O[100:36], IN1);
  UBZero_35_35 U2 (O[35]);
  UB1DCON_34 U3 (O[34], IN2);
endmodule

module UBCMBIN_103_103_1000 (O, IN0, IN1, IN2);
  output [103:36] O;
  input IN0;
  input [102:38] IN1;
  input IN2;
  UB1DCON_103 U0 (O[103], IN0);
  UBCON_102_38 U1 (O[102:38], IN1);
  UBZero_37_37 U2 (O[37]);
  UB1DCON_36 U3 (O[36], IN2);
endmodule

module UBCMBIN_105_105_1000 (O, IN0, IN1, IN2);
  output [105:38] O;
  input IN0;
  input [104:40] IN1;
  input IN2;
  UB1DCON_105 U0 (O[105], IN0);
  UBCON_104_40 U1 (O[104:40], IN1);
  UBZero_39_39 U2 (O[39]);
  UB1DCON_38 U3 (O[38], IN2);
endmodule

module UBCMBIN_107_107_1000 (O, IN0, IN1, IN2);
  output [107:40] O;
  input IN0;
  input [106:42] IN1;
  input IN2;
  UB1DCON_107 U0 (O[107], IN0);
  UBCON_106_42 U1 (O[106:42], IN1);
  UBZero_41_41 U2 (O[41]);
  UB1DCON_40 U3 (O[40], IN2);
endmodule

module UBCMBIN_109_109_1000 (O, IN0, IN1, IN2);
  output [109:42] O;
  input IN0;
  input [108:44] IN1;
  input IN2;
  UB1DCON_109 U0 (O[109], IN0);
  UBCON_108_44 U1 (O[108:44], IN1);
  UBZero_43_43 U2 (O[43]);
  UB1DCON_42 U3 (O[42], IN2);
endmodule

module UBCMBIN_111_111_1000 (O, IN0, IN1, IN2);
  output [111:44] O;
  input IN0;
  input [110:46] IN1;
  input IN2;
  UB1DCON_111 U0 (O[111], IN0);
  UBCON_110_46 U1 (O[110:46], IN1);
  UBZero_45_45 U2 (O[45]);
  UB1DCON_44 U3 (O[44], IN2);
endmodule

module UBCMBIN_113_113_1000 (O, IN0, IN1, IN2);
  output [113:46] O;
  input IN0;
  input [112:48] IN1;
  input IN2;
  UB1DCON_113 U0 (O[113], IN0);
  UBCON_112_48 U1 (O[112:48], IN1);
  UBZero_47_47 U2 (O[47]);
  UB1DCON_46 U3 (O[46], IN2);
endmodule

module UBCMBIN_115_115_1000 (O, IN0, IN1, IN2);
  output [115:48] O;
  input IN0;
  input [114:50] IN1;
  input IN2;
  UB1DCON_115 U0 (O[115], IN0);
  UBCON_114_50 U1 (O[114:50], IN1);
  UBZero_49_49 U2 (O[49]);
  UB1DCON_48 U3 (O[48], IN2);
endmodule

module UBCMBIN_117_117_1000 (O, IN0, IN1, IN2);
  output [117:50] O;
  input IN0;
  input [116:52] IN1;
  input IN2;
  UB1DCON_117 U0 (O[117], IN0);
  UBCON_116_52 U1 (O[116:52], IN1);
  UBZero_51_51 U2 (O[51]);
  UB1DCON_50 U3 (O[50], IN2);
endmodule

module UBCMBIN_119_119_1000 (O, IN0, IN1, IN2);
  output [119:52] O;
  input IN0;
  input [118:54] IN1;
  input IN2;
  UB1DCON_119 U0 (O[119], IN0);
  UBCON_118_54 U1 (O[118:54], IN1);
  UBZero_53_53 U2 (O[53]);
  UB1DCON_52 U3 (O[52], IN2);
endmodule

module UBCMBIN_121_121_1000 (O, IN0, IN1, IN2);
  output [121:54] O;
  input IN0;
  input [120:56] IN1;
  input IN2;
  UB1DCON_121 U0 (O[121], IN0);
  UBCON_120_56 U1 (O[120:56], IN1);
  UBZero_55_55 U2 (O[55]);
  UB1DCON_54 U3 (O[54], IN2);
endmodule

module UBCMBIN_123_123_1000 (O, IN0, IN1, IN2);
  output [123:56] O;
  input IN0;
  input [122:58] IN1;
  input IN2;
  UB1DCON_123 U0 (O[123], IN0);
  UBCON_122_58 U1 (O[122:58], IN1);
  UBZero_57_57 U2 (O[57]);
  UB1DCON_56 U3 (O[56], IN2);
endmodule

module UBCMBIN_125_125_1000 (O, IN0, IN1, IN2);
  output [125:58] O;
  input IN0;
  input [124:60] IN1;
  input IN2;
  UB1DCON_125 U0 (O[125], IN0);
  UBCON_124_60 U1 (O[124:60], IN1);
  UBZero_59_59 U2 (O[59]);
  UB1DCON_58 U3 (O[58], IN2);
endmodule

module UBCMBIN_126_62_60000 (O, IN0, IN1);
  output [126:60] O;
  input [126:62] IN0;
  input IN1;
  UBCON_126_62 U0 (O[126:62], IN0);
  UBZero_61_61 U1 (O[61]);
  UB1DCON_60 U2 (O[60], IN1);
endmodule

module UBCMBIN_64_64_62_000 (O, IN0, IN1);
  output [64:62] O;
  input IN0;
  input IN1;
  UB1DCON_64 U0 (O[64], IN0);
  UBZero_63_63 U1 (O[63]);
  UB1DCON_62 U2 (O[62], IN1);
endmodule

module UBCMBIN_65_65_64_000 (O, IN0, IN1);
  output [65:0] O;
  input IN0;
  input [64:0] IN1;
  UB1DCON_65 U0 (O[65], IN0);
  UBCON_64_0 U1 (O[64:0], IN1);
endmodule

module UBCMBIN_67_67_66_000 (O, IN0, IN1, IN2);
  output [67:0] O;
  input IN0;
  input [66:2] IN1;
  input IN2;
  UB1DCON_67 U0 (O[67], IN0);
  UBCON_66_2 U1 (O[66:2], IN1);
  UBZero_1_1 U2 (O[1]);
  UB1DCON_0 U3 (O[0], IN2);
endmodule

module UBCMBIN_69_69_68_000 (O, IN0, IN1, IN2);
  output [69:2] O;
  input IN0;
  input [68:4] IN1;
  input IN2;
  UB1DCON_69 U0 (O[69], IN0);
  UBCON_68_4 U1 (O[68:4], IN1);
  UBZero_3_3 U2 (O[3]);
  UB1DCON_2 U3 (O[2], IN2);
endmodule

module UBCMBIN_71_71_70_000 (O, IN0, IN1, IN2);
  output [71:4] O;
  input IN0;
  input [70:6] IN1;
  input IN2;
  UB1DCON_71 U0 (O[71], IN0);
  UBCON_70_6 U1 (O[70:6], IN1);
  UBZero_5_5 U2 (O[5]);
  UB1DCON_4 U3 (O[4], IN2);
endmodule

module UBCMBIN_73_73_72_000 (O, IN0, IN1, IN2);
  output [73:6] O;
  input IN0;
  input [72:8] IN1;
  input IN2;
  UB1DCON_73 U0 (O[73], IN0);
  UBCON_72_8 U1 (O[72:8], IN1);
  UBZero_7_7 U2 (O[7]);
  UB1DCON_6 U3 (O[6], IN2);
endmodule

module UBCMBIN_75_75_74_000 (O, IN0, IN1, IN2);
  output [75:8] O;
  input IN0;
  input [74:10] IN1;
  input IN2;
  UB1DCON_75 U0 (O[75], IN0);
  UBCON_74_10 U1 (O[74:10], IN1);
  UBZero_9_9 U2 (O[9]);
  UB1DCON_8 U3 (O[8], IN2);
endmodule

module UBCMBIN_77_77_76_000 (O, IN0, IN1, IN2);
  output [77:10] O;
  input IN0;
  input [76:12] IN1;
  input IN2;
  UB1DCON_77 U0 (O[77], IN0);
  UBCON_76_12 U1 (O[76:12], IN1);
  UBZero_11_11 U2 (O[11]);
  UB1DCON_10 U3 (O[10], IN2);
endmodule

module UBCMBIN_79_79_78_000 (O, IN0, IN1, IN2);
  output [79:12] O;
  input IN0;
  input [78:14] IN1;
  input IN2;
  UB1DCON_79 U0 (O[79], IN0);
  UBCON_78_14 U1 (O[78:14], IN1);
  UBZero_13_13 U2 (O[13]);
  UB1DCON_12 U3 (O[12], IN2);
endmodule

module UBCMBIN_81_81_80_000 (O, IN0, IN1, IN2);
  output [81:14] O;
  input IN0;
  input [80:16] IN1;
  input IN2;
  UB1DCON_81 U0 (O[81], IN0);
  UBCON_80_16 U1 (O[80:16], IN1);
  UBZero_15_15 U2 (O[15]);
  UB1DCON_14 U3 (O[14], IN2);
endmodule

module UBCMBIN_83_83_82_000 (O, IN0, IN1, IN2);
  output [83:16] O;
  input IN0;
  input [82:18] IN1;
  input IN2;
  UB1DCON_83 U0 (O[83], IN0);
  UBCON_82_18 U1 (O[82:18], IN1);
  UBZero_17_17 U2 (O[17]);
  UB1DCON_16 U3 (O[16], IN2);
endmodule

module UBCMBIN_85_85_84_000 (O, IN0, IN1, IN2);
  output [85:18] O;
  input IN0;
  input [84:20] IN1;
  input IN2;
  UB1DCON_85 U0 (O[85], IN0);
  UBCON_84_20 U1 (O[84:20], IN1);
  UBZero_19_19 U2 (O[19]);
  UB1DCON_18 U3 (O[18], IN2);
endmodule

module UBCMBIN_87_87_86_000 (O, IN0, IN1, IN2);
  output [87:20] O;
  input IN0;
  input [86:22] IN1;
  input IN2;
  UB1DCON_87 U0 (O[87], IN0);
  UBCON_86_22 U1 (O[86:22], IN1);
  UBZero_21_21 U2 (O[21]);
  UB1DCON_20 U3 (O[20], IN2);
endmodule

module UBCMBIN_89_89_88_000 (O, IN0, IN1, IN2);
  output [89:22] O;
  input IN0;
  input [88:24] IN1;
  input IN2;
  UB1DCON_89 U0 (O[89], IN0);
  UBCON_88_24 U1 (O[88:24], IN1);
  UBZero_23_23 U2 (O[23]);
  UB1DCON_22 U3 (O[22], IN2);
endmodule

module UBCMBIN_91_91_90_000 (O, IN0, IN1, IN2);
  output [91:24] O;
  input IN0;
  input [90:26] IN1;
  input IN2;
  UB1DCON_91 U0 (O[91], IN0);
  UBCON_90_26 U1 (O[90:26], IN1);
  UBZero_25_25 U2 (O[25]);
  UB1DCON_24 U3 (O[24], IN2);
endmodule

module UBCMBIN_93_93_92_000 (O, IN0, IN1, IN2);
  output [93:26] O;
  input IN0;
  input [92:28] IN1;
  input IN2;
  UB1DCON_93 U0 (O[93], IN0);
  UBCON_92_28 U1 (O[92:28], IN1);
  UBZero_27_27 U2 (O[27]);
  UB1DCON_26 U3 (O[26], IN2);
endmodule

module UBCMBIN_95_95_94_000 (O, IN0, IN1, IN2);
  output [95:28] O;
  input IN0;
  input [94:30] IN1;
  input IN2;
  UB1DCON_95 U0 (O[95], IN0);
  UBCON_94_30 U1 (O[94:30], IN1);
  UBZero_29_29 U2 (O[29]);
  UB1DCON_28 U3 (O[28], IN2);
endmodule

module UBCMBIN_97_97_96_000 (O, IN0, IN1, IN2);
  output [97:30] O;
  input IN0;
  input [96:32] IN1;
  input IN2;
  UB1DCON_97 U0 (O[97], IN0);
  UBCON_96_32 U1 (O[96:32], IN1);
  UBZero_31_31 U2 (O[31]);
  UB1DCON_30 U3 (O[30], IN2);
endmodule

module UBCMBIN_99_99_98_000 (O, IN0, IN1, IN2);
  output [99:32] O;
  input IN0;
  input [98:34] IN1;
  input IN2;
  UB1DCON_99 U0 (O[99], IN0);
  UBCON_98_34 U1 (O[98:34], IN1);
  UBZero_33_33 U2 (O[33]);
  UB1DCON_32 U3 (O[32], IN2);
endmodule

module UBCON_100_26 (O, I);
  output [100:26] O;
  input [100:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
  UB1DCON_28 U2 (O[28], I[28]);
  UB1DCON_29 U3 (O[29], I[29]);
  UB1DCON_30 U4 (O[30], I[30]);
  UB1DCON_31 U5 (O[31], I[31]);
  UB1DCON_32 U6 (O[32], I[32]);
  UB1DCON_33 U7 (O[33], I[33]);
  UB1DCON_34 U8 (O[34], I[34]);
  UB1DCON_35 U9 (O[35], I[35]);
  UB1DCON_36 U10 (O[36], I[36]);
  UB1DCON_37 U11 (O[37], I[37]);
  UB1DCON_38 U12 (O[38], I[38]);
  UB1DCON_39 U13 (O[39], I[39]);
  UB1DCON_40 U14 (O[40], I[40]);
  UB1DCON_41 U15 (O[41], I[41]);
  UB1DCON_42 U16 (O[42], I[42]);
  UB1DCON_43 U17 (O[43], I[43]);
  UB1DCON_44 U18 (O[44], I[44]);
  UB1DCON_45 U19 (O[45], I[45]);
  UB1DCON_46 U20 (O[46], I[46]);
  UB1DCON_47 U21 (O[47], I[47]);
  UB1DCON_48 U22 (O[48], I[48]);
  UB1DCON_49 U23 (O[49], I[49]);
  UB1DCON_50 U24 (O[50], I[50]);
  UB1DCON_51 U25 (O[51], I[51]);
  UB1DCON_52 U26 (O[52], I[52]);
  UB1DCON_53 U27 (O[53], I[53]);
  UB1DCON_54 U28 (O[54], I[54]);
  UB1DCON_55 U29 (O[55], I[55]);
  UB1DCON_56 U30 (O[56], I[56]);
  UB1DCON_57 U31 (O[57], I[57]);
  UB1DCON_58 U32 (O[58], I[58]);
  UB1DCON_59 U33 (O[59], I[59]);
  UB1DCON_60 U34 (O[60], I[60]);
  UB1DCON_61 U35 (O[61], I[61]);
  UB1DCON_62 U36 (O[62], I[62]);
  UB1DCON_63 U37 (O[63], I[63]);
  UB1DCON_64 U38 (O[64], I[64]);
  UB1DCON_65 U39 (O[65], I[65]);
  UB1DCON_66 U40 (O[66], I[66]);
  UB1DCON_67 U41 (O[67], I[67]);
  UB1DCON_68 U42 (O[68], I[68]);
  UB1DCON_69 U43 (O[69], I[69]);
  UB1DCON_70 U44 (O[70], I[70]);
  UB1DCON_71 U45 (O[71], I[71]);
  UB1DCON_72 U46 (O[72], I[72]);
  UB1DCON_73 U47 (O[73], I[73]);
  UB1DCON_74 U48 (O[74], I[74]);
  UB1DCON_75 U49 (O[75], I[75]);
  UB1DCON_76 U50 (O[76], I[76]);
  UB1DCON_77 U51 (O[77], I[77]);
  UB1DCON_78 U52 (O[78], I[78]);
  UB1DCON_79 U53 (O[79], I[79]);
  UB1DCON_80 U54 (O[80], I[80]);
  UB1DCON_81 U55 (O[81], I[81]);
  UB1DCON_82 U56 (O[82], I[82]);
  UB1DCON_83 U57 (O[83], I[83]);
  UB1DCON_84 U58 (O[84], I[84]);
  UB1DCON_85 U59 (O[85], I[85]);
  UB1DCON_86 U60 (O[86], I[86]);
  UB1DCON_87 U61 (O[87], I[87]);
  UB1DCON_88 U62 (O[88], I[88]);
  UB1DCON_89 U63 (O[89], I[89]);
  UB1DCON_90 U64 (O[90], I[90]);
  UB1DCON_91 U65 (O[91], I[91]);
  UB1DCON_92 U66 (O[92], I[92]);
  UB1DCON_93 U67 (O[93], I[93]);
  UB1DCON_94 U68 (O[94], I[94]);
  UB1DCON_95 U69 (O[95], I[95]);
  UB1DCON_96 U70 (O[96], I[96]);
  UB1DCON_97 U71 (O[97], I[97]);
  UB1DCON_98 U72 (O[98], I[98]);
  UB1DCON_99 U73 (O[99], I[99]);
  UB1DCON_100 U74 (O[100], I[100]);
endmodule

module UBCON_100_36 (O, I);
  output [100:36] O;
  input [100:36] I;
  UB1DCON_36 U0 (O[36], I[36]);
  UB1DCON_37 U1 (O[37], I[37]);
  UB1DCON_38 U2 (O[38], I[38]);
  UB1DCON_39 U3 (O[39], I[39]);
  UB1DCON_40 U4 (O[40], I[40]);
  UB1DCON_41 U5 (O[41], I[41]);
  UB1DCON_42 U6 (O[42], I[42]);
  UB1DCON_43 U7 (O[43], I[43]);
  UB1DCON_44 U8 (O[44], I[44]);
  UB1DCON_45 U9 (O[45], I[45]);
  UB1DCON_46 U10 (O[46], I[46]);
  UB1DCON_47 U11 (O[47], I[47]);
  UB1DCON_48 U12 (O[48], I[48]);
  UB1DCON_49 U13 (O[49], I[49]);
  UB1DCON_50 U14 (O[50], I[50]);
  UB1DCON_51 U15 (O[51], I[51]);
  UB1DCON_52 U16 (O[52], I[52]);
  UB1DCON_53 U17 (O[53], I[53]);
  UB1DCON_54 U18 (O[54], I[54]);
  UB1DCON_55 U19 (O[55], I[55]);
  UB1DCON_56 U20 (O[56], I[56]);
  UB1DCON_57 U21 (O[57], I[57]);
  UB1DCON_58 U22 (O[58], I[58]);
  UB1DCON_59 U23 (O[59], I[59]);
  UB1DCON_60 U24 (O[60], I[60]);
  UB1DCON_61 U25 (O[61], I[61]);
  UB1DCON_62 U26 (O[62], I[62]);
  UB1DCON_63 U27 (O[63], I[63]);
  UB1DCON_64 U28 (O[64], I[64]);
  UB1DCON_65 U29 (O[65], I[65]);
  UB1DCON_66 U30 (O[66], I[66]);
  UB1DCON_67 U31 (O[67], I[67]);
  UB1DCON_68 U32 (O[68], I[68]);
  UB1DCON_69 U33 (O[69], I[69]);
  UB1DCON_70 U34 (O[70], I[70]);
  UB1DCON_71 U35 (O[71], I[71]);
  UB1DCON_72 U36 (O[72], I[72]);
  UB1DCON_73 U37 (O[73], I[73]);
  UB1DCON_74 U38 (O[74], I[74]);
  UB1DCON_75 U39 (O[75], I[75]);
  UB1DCON_76 U40 (O[76], I[76]);
  UB1DCON_77 U41 (O[77], I[77]);
  UB1DCON_78 U42 (O[78], I[78]);
  UB1DCON_79 U43 (O[79], I[79]);
  UB1DCON_80 U44 (O[80], I[80]);
  UB1DCON_81 U45 (O[81], I[81]);
  UB1DCON_82 U46 (O[82], I[82]);
  UB1DCON_83 U47 (O[83], I[83]);
  UB1DCON_84 U48 (O[84], I[84]);
  UB1DCON_85 U49 (O[85], I[85]);
  UB1DCON_86 U50 (O[86], I[86]);
  UB1DCON_87 U51 (O[87], I[87]);
  UB1DCON_88 U52 (O[88], I[88]);
  UB1DCON_89 U53 (O[89], I[89]);
  UB1DCON_90 U54 (O[90], I[90]);
  UB1DCON_91 U55 (O[91], I[91]);
  UB1DCON_92 U56 (O[92], I[92]);
  UB1DCON_93 U57 (O[93], I[93]);
  UB1DCON_94 U58 (O[94], I[94]);
  UB1DCON_95 U59 (O[95], I[95]);
  UB1DCON_96 U60 (O[96], I[96]);
  UB1DCON_97 U61 (O[97], I[97]);
  UB1DCON_98 U62 (O[98], I[98]);
  UB1DCON_99 U63 (O[99], I[99]);
  UB1DCON_100 U64 (O[100], I[100]);
endmodule

module UBCON_101_100 (O, I);
  output [101:100] O;
  input [101:100] I;
  UB1DCON_100 U0 (O[100], I[100]);
  UB1DCON_101 U1 (O[101], I[101]);
endmodule

module UBCON_102_38 (O, I);
  output [102:38] O;
  input [102:38] I;
  UB1DCON_38 U0 (O[38], I[38]);
  UB1DCON_39 U1 (O[39], I[39]);
  UB1DCON_40 U2 (O[40], I[40]);
  UB1DCON_41 U3 (O[41], I[41]);
  UB1DCON_42 U4 (O[42], I[42]);
  UB1DCON_43 U5 (O[43], I[43]);
  UB1DCON_44 U6 (O[44], I[44]);
  UB1DCON_45 U7 (O[45], I[45]);
  UB1DCON_46 U8 (O[46], I[46]);
  UB1DCON_47 U9 (O[47], I[47]);
  UB1DCON_48 U10 (O[48], I[48]);
  UB1DCON_49 U11 (O[49], I[49]);
  UB1DCON_50 U12 (O[50], I[50]);
  UB1DCON_51 U13 (O[51], I[51]);
  UB1DCON_52 U14 (O[52], I[52]);
  UB1DCON_53 U15 (O[53], I[53]);
  UB1DCON_54 U16 (O[54], I[54]);
  UB1DCON_55 U17 (O[55], I[55]);
  UB1DCON_56 U18 (O[56], I[56]);
  UB1DCON_57 U19 (O[57], I[57]);
  UB1DCON_58 U20 (O[58], I[58]);
  UB1DCON_59 U21 (O[59], I[59]);
  UB1DCON_60 U22 (O[60], I[60]);
  UB1DCON_61 U23 (O[61], I[61]);
  UB1DCON_62 U24 (O[62], I[62]);
  UB1DCON_63 U25 (O[63], I[63]);
  UB1DCON_64 U26 (O[64], I[64]);
  UB1DCON_65 U27 (O[65], I[65]);
  UB1DCON_66 U28 (O[66], I[66]);
  UB1DCON_67 U29 (O[67], I[67]);
  UB1DCON_68 U30 (O[68], I[68]);
  UB1DCON_69 U31 (O[69], I[69]);
  UB1DCON_70 U32 (O[70], I[70]);
  UB1DCON_71 U33 (O[71], I[71]);
  UB1DCON_72 U34 (O[72], I[72]);
  UB1DCON_73 U35 (O[73], I[73]);
  UB1DCON_74 U36 (O[74], I[74]);
  UB1DCON_75 U37 (O[75], I[75]);
  UB1DCON_76 U38 (O[76], I[76]);
  UB1DCON_77 U39 (O[77], I[77]);
  UB1DCON_78 U40 (O[78], I[78]);
  UB1DCON_79 U41 (O[79], I[79]);
  UB1DCON_80 U42 (O[80], I[80]);
  UB1DCON_81 U43 (O[81], I[81]);
  UB1DCON_82 U44 (O[82], I[82]);
  UB1DCON_83 U45 (O[83], I[83]);
  UB1DCON_84 U46 (O[84], I[84]);
  UB1DCON_85 U47 (O[85], I[85]);
  UB1DCON_86 U48 (O[86], I[86]);
  UB1DCON_87 U49 (O[87], I[87]);
  UB1DCON_88 U50 (O[88], I[88]);
  UB1DCON_89 U51 (O[89], I[89]);
  UB1DCON_90 U52 (O[90], I[90]);
  UB1DCON_91 U53 (O[91], I[91]);
  UB1DCON_92 U54 (O[92], I[92]);
  UB1DCON_93 U55 (O[93], I[93]);
  UB1DCON_94 U56 (O[94], I[94]);
  UB1DCON_95 U57 (O[95], I[95]);
  UB1DCON_96 U58 (O[96], I[96]);
  UB1DCON_97 U59 (O[97], I[97]);
  UB1DCON_98 U60 (O[98], I[98]);
  UB1DCON_99 U61 (O[99], I[99]);
  UB1DCON_100 U62 (O[100], I[100]);
  UB1DCON_101 U63 (O[101], I[101]);
  UB1DCON_102 U64 (O[102], I[102]);
endmodule

module UBCON_103_102 (O, I);
  output [103:102] O;
  input [103:102] I;
  UB1DCON_102 U0 (O[102], I[102]);
  UB1DCON_103 U1 (O[103], I[103]);
endmodule

module UBCON_104_40 (O, I);
  output [104:40] O;
  input [104:40] I;
  UB1DCON_40 U0 (O[40], I[40]);
  UB1DCON_41 U1 (O[41], I[41]);
  UB1DCON_42 U2 (O[42], I[42]);
  UB1DCON_43 U3 (O[43], I[43]);
  UB1DCON_44 U4 (O[44], I[44]);
  UB1DCON_45 U5 (O[45], I[45]);
  UB1DCON_46 U6 (O[46], I[46]);
  UB1DCON_47 U7 (O[47], I[47]);
  UB1DCON_48 U8 (O[48], I[48]);
  UB1DCON_49 U9 (O[49], I[49]);
  UB1DCON_50 U10 (O[50], I[50]);
  UB1DCON_51 U11 (O[51], I[51]);
  UB1DCON_52 U12 (O[52], I[52]);
  UB1DCON_53 U13 (O[53], I[53]);
  UB1DCON_54 U14 (O[54], I[54]);
  UB1DCON_55 U15 (O[55], I[55]);
  UB1DCON_56 U16 (O[56], I[56]);
  UB1DCON_57 U17 (O[57], I[57]);
  UB1DCON_58 U18 (O[58], I[58]);
  UB1DCON_59 U19 (O[59], I[59]);
  UB1DCON_60 U20 (O[60], I[60]);
  UB1DCON_61 U21 (O[61], I[61]);
  UB1DCON_62 U22 (O[62], I[62]);
  UB1DCON_63 U23 (O[63], I[63]);
  UB1DCON_64 U24 (O[64], I[64]);
  UB1DCON_65 U25 (O[65], I[65]);
  UB1DCON_66 U26 (O[66], I[66]);
  UB1DCON_67 U27 (O[67], I[67]);
  UB1DCON_68 U28 (O[68], I[68]);
  UB1DCON_69 U29 (O[69], I[69]);
  UB1DCON_70 U30 (O[70], I[70]);
  UB1DCON_71 U31 (O[71], I[71]);
  UB1DCON_72 U32 (O[72], I[72]);
  UB1DCON_73 U33 (O[73], I[73]);
  UB1DCON_74 U34 (O[74], I[74]);
  UB1DCON_75 U35 (O[75], I[75]);
  UB1DCON_76 U36 (O[76], I[76]);
  UB1DCON_77 U37 (O[77], I[77]);
  UB1DCON_78 U38 (O[78], I[78]);
  UB1DCON_79 U39 (O[79], I[79]);
  UB1DCON_80 U40 (O[80], I[80]);
  UB1DCON_81 U41 (O[81], I[81]);
  UB1DCON_82 U42 (O[82], I[82]);
  UB1DCON_83 U43 (O[83], I[83]);
  UB1DCON_84 U44 (O[84], I[84]);
  UB1DCON_85 U45 (O[85], I[85]);
  UB1DCON_86 U46 (O[86], I[86]);
  UB1DCON_87 U47 (O[87], I[87]);
  UB1DCON_88 U48 (O[88], I[88]);
  UB1DCON_89 U49 (O[89], I[89]);
  UB1DCON_90 U50 (O[90], I[90]);
  UB1DCON_91 U51 (O[91], I[91]);
  UB1DCON_92 U52 (O[92], I[92]);
  UB1DCON_93 U53 (O[93], I[93]);
  UB1DCON_94 U54 (O[94], I[94]);
  UB1DCON_95 U55 (O[95], I[95]);
  UB1DCON_96 U56 (O[96], I[96]);
  UB1DCON_97 U57 (O[97], I[97]);
  UB1DCON_98 U58 (O[98], I[98]);
  UB1DCON_99 U59 (O[99], I[99]);
  UB1DCON_100 U60 (O[100], I[100]);
  UB1DCON_101 U61 (O[101], I[101]);
  UB1DCON_102 U62 (O[102], I[102]);
  UB1DCON_103 U63 (O[103], I[103]);
  UB1DCON_104 U64 (O[104], I[104]);
endmodule

module UBCON_105_104 (O, I);
  output [105:104] O;
  input [105:104] I;
  UB1DCON_104 U0 (O[104], I[104]);
  UB1DCON_105 U1 (O[105], I[105]);
endmodule

module UBCON_106_42 (O, I);
  output [106:42] O;
  input [106:42] I;
  UB1DCON_42 U0 (O[42], I[42]);
  UB1DCON_43 U1 (O[43], I[43]);
  UB1DCON_44 U2 (O[44], I[44]);
  UB1DCON_45 U3 (O[45], I[45]);
  UB1DCON_46 U4 (O[46], I[46]);
  UB1DCON_47 U5 (O[47], I[47]);
  UB1DCON_48 U6 (O[48], I[48]);
  UB1DCON_49 U7 (O[49], I[49]);
  UB1DCON_50 U8 (O[50], I[50]);
  UB1DCON_51 U9 (O[51], I[51]);
  UB1DCON_52 U10 (O[52], I[52]);
  UB1DCON_53 U11 (O[53], I[53]);
  UB1DCON_54 U12 (O[54], I[54]);
  UB1DCON_55 U13 (O[55], I[55]);
  UB1DCON_56 U14 (O[56], I[56]);
  UB1DCON_57 U15 (O[57], I[57]);
  UB1DCON_58 U16 (O[58], I[58]);
  UB1DCON_59 U17 (O[59], I[59]);
  UB1DCON_60 U18 (O[60], I[60]);
  UB1DCON_61 U19 (O[61], I[61]);
  UB1DCON_62 U20 (O[62], I[62]);
  UB1DCON_63 U21 (O[63], I[63]);
  UB1DCON_64 U22 (O[64], I[64]);
  UB1DCON_65 U23 (O[65], I[65]);
  UB1DCON_66 U24 (O[66], I[66]);
  UB1DCON_67 U25 (O[67], I[67]);
  UB1DCON_68 U26 (O[68], I[68]);
  UB1DCON_69 U27 (O[69], I[69]);
  UB1DCON_70 U28 (O[70], I[70]);
  UB1DCON_71 U29 (O[71], I[71]);
  UB1DCON_72 U30 (O[72], I[72]);
  UB1DCON_73 U31 (O[73], I[73]);
  UB1DCON_74 U32 (O[74], I[74]);
  UB1DCON_75 U33 (O[75], I[75]);
  UB1DCON_76 U34 (O[76], I[76]);
  UB1DCON_77 U35 (O[77], I[77]);
  UB1DCON_78 U36 (O[78], I[78]);
  UB1DCON_79 U37 (O[79], I[79]);
  UB1DCON_80 U38 (O[80], I[80]);
  UB1DCON_81 U39 (O[81], I[81]);
  UB1DCON_82 U40 (O[82], I[82]);
  UB1DCON_83 U41 (O[83], I[83]);
  UB1DCON_84 U42 (O[84], I[84]);
  UB1DCON_85 U43 (O[85], I[85]);
  UB1DCON_86 U44 (O[86], I[86]);
  UB1DCON_87 U45 (O[87], I[87]);
  UB1DCON_88 U46 (O[88], I[88]);
  UB1DCON_89 U47 (O[89], I[89]);
  UB1DCON_90 U48 (O[90], I[90]);
  UB1DCON_91 U49 (O[91], I[91]);
  UB1DCON_92 U50 (O[92], I[92]);
  UB1DCON_93 U51 (O[93], I[93]);
  UB1DCON_94 U52 (O[94], I[94]);
  UB1DCON_95 U53 (O[95], I[95]);
  UB1DCON_96 U54 (O[96], I[96]);
  UB1DCON_97 U55 (O[97], I[97]);
  UB1DCON_98 U56 (O[98], I[98]);
  UB1DCON_99 U57 (O[99], I[99]);
  UB1DCON_100 U58 (O[100], I[100]);
  UB1DCON_101 U59 (O[101], I[101]);
  UB1DCON_102 U60 (O[102], I[102]);
  UB1DCON_103 U61 (O[103], I[103]);
  UB1DCON_104 U62 (O[104], I[104]);
  UB1DCON_105 U63 (O[105], I[105]);
  UB1DCON_106 U64 (O[106], I[106]);
endmodule

module UBCON_107_106 (O, I);
  output [107:106] O;
  input [107:106] I;
  UB1DCON_106 U0 (O[106], I[106]);
  UB1DCON_107 U1 (O[107], I[107]);
endmodule

module UBCON_108_44 (O, I);
  output [108:44] O;
  input [108:44] I;
  UB1DCON_44 U0 (O[44], I[44]);
  UB1DCON_45 U1 (O[45], I[45]);
  UB1DCON_46 U2 (O[46], I[46]);
  UB1DCON_47 U3 (O[47], I[47]);
  UB1DCON_48 U4 (O[48], I[48]);
  UB1DCON_49 U5 (O[49], I[49]);
  UB1DCON_50 U6 (O[50], I[50]);
  UB1DCON_51 U7 (O[51], I[51]);
  UB1DCON_52 U8 (O[52], I[52]);
  UB1DCON_53 U9 (O[53], I[53]);
  UB1DCON_54 U10 (O[54], I[54]);
  UB1DCON_55 U11 (O[55], I[55]);
  UB1DCON_56 U12 (O[56], I[56]);
  UB1DCON_57 U13 (O[57], I[57]);
  UB1DCON_58 U14 (O[58], I[58]);
  UB1DCON_59 U15 (O[59], I[59]);
  UB1DCON_60 U16 (O[60], I[60]);
  UB1DCON_61 U17 (O[61], I[61]);
  UB1DCON_62 U18 (O[62], I[62]);
  UB1DCON_63 U19 (O[63], I[63]);
  UB1DCON_64 U20 (O[64], I[64]);
  UB1DCON_65 U21 (O[65], I[65]);
  UB1DCON_66 U22 (O[66], I[66]);
  UB1DCON_67 U23 (O[67], I[67]);
  UB1DCON_68 U24 (O[68], I[68]);
  UB1DCON_69 U25 (O[69], I[69]);
  UB1DCON_70 U26 (O[70], I[70]);
  UB1DCON_71 U27 (O[71], I[71]);
  UB1DCON_72 U28 (O[72], I[72]);
  UB1DCON_73 U29 (O[73], I[73]);
  UB1DCON_74 U30 (O[74], I[74]);
  UB1DCON_75 U31 (O[75], I[75]);
  UB1DCON_76 U32 (O[76], I[76]);
  UB1DCON_77 U33 (O[77], I[77]);
  UB1DCON_78 U34 (O[78], I[78]);
  UB1DCON_79 U35 (O[79], I[79]);
  UB1DCON_80 U36 (O[80], I[80]);
  UB1DCON_81 U37 (O[81], I[81]);
  UB1DCON_82 U38 (O[82], I[82]);
  UB1DCON_83 U39 (O[83], I[83]);
  UB1DCON_84 U40 (O[84], I[84]);
  UB1DCON_85 U41 (O[85], I[85]);
  UB1DCON_86 U42 (O[86], I[86]);
  UB1DCON_87 U43 (O[87], I[87]);
  UB1DCON_88 U44 (O[88], I[88]);
  UB1DCON_89 U45 (O[89], I[89]);
  UB1DCON_90 U46 (O[90], I[90]);
  UB1DCON_91 U47 (O[91], I[91]);
  UB1DCON_92 U48 (O[92], I[92]);
  UB1DCON_93 U49 (O[93], I[93]);
  UB1DCON_94 U50 (O[94], I[94]);
  UB1DCON_95 U51 (O[95], I[95]);
  UB1DCON_96 U52 (O[96], I[96]);
  UB1DCON_97 U53 (O[97], I[97]);
  UB1DCON_98 U54 (O[98], I[98]);
  UB1DCON_99 U55 (O[99], I[99]);
  UB1DCON_100 U56 (O[100], I[100]);
  UB1DCON_101 U57 (O[101], I[101]);
  UB1DCON_102 U58 (O[102], I[102]);
  UB1DCON_103 U59 (O[103], I[103]);
  UB1DCON_104 U60 (O[104], I[104]);
  UB1DCON_105 U61 (O[105], I[105]);
  UB1DCON_106 U62 (O[106], I[106]);
  UB1DCON_107 U63 (O[107], I[107]);
  UB1DCON_108 U64 (O[108], I[108]);
endmodule

module UBCON_109_108 (O, I);
  output [109:108] O;
  input [109:108] I;
  UB1DCON_108 U0 (O[108], I[108]);
  UB1DCON_109 U1 (O[109], I[109]);
endmodule

module UBCON_110_46 (O, I);
  output [110:46] O;
  input [110:46] I;
  UB1DCON_46 U0 (O[46], I[46]);
  UB1DCON_47 U1 (O[47], I[47]);
  UB1DCON_48 U2 (O[48], I[48]);
  UB1DCON_49 U3 (O[49], I[49]);
  UB1DCON_50 U4 (O[50], I[50]);
  UB1DCON_51 U5 (O[51], I[51]);
  UB1DCON_52 U6 (O[52], I[52]);
  UB1DCON_53 U7 (O[53], I[53]);
  UB1DCON_54 U8 (O[54], I[54]);
  UB1DCON_55 U9 (O[55], I[55]);
  UB1DCON_56 U10 (O[56], I[56]);
  UB1DCON_57 U11 (O[57], I[57]);
  UB1DCON_58 U12 (O[58], I[58]);
  UB1DCON_59 U13 (O[59], I[59]);
  UB1DCON_60 U14 (O[60], I[60]);
  UB1DCON_61 U15 (O[61], I[61]);
  UB1DCON_62 U16 (O[62], I[62]);
  UB1DCON_63 U17 (O[63], I[63]);
  UB1DCON_64 U18 (O[64], I[64]);
  UB1DCON_65 U19 (O[65], I[65]);
  UB1DCON_66 U20 (O[66], I[66]);
  UB1DCON_67 U21 (O[67], I[67]);
  UB1DCON_68 U22 (O[68], I[68]);
  UB1DCON_69 U23 (O[69], I[69]);
  UB1DCON_70 U24 (O[70], I[70]);
  UB1DCON_71 U25 (O[71], I[71]);
  UB1DCON_72 U26 (O[72], I[72]);
  UB1DCON_73 U27 (O[73], I[73]);
  UB1DCON_74 U28 (O[74], I[74]);
  UB1DCON_75 U29 (O[75], I[75]);
  UB1DCON_76 U30 (O[76], I[76]);
  UB1DCON_77 U31 (O[77], I[77]);
  UB1DCON_78 U32 (O[78], I[78]);
  UB1DCON_79 U33 (O[79], I[79]);
  UB1DCON_80 U34 (O[80], I[80]);
  UB1DCON_81 U35 (O[81], I[81]);
  UB1DCON_82 U36 (O[82], I[82]);
  UB1DCON_83 U37 (O[83], I[83]);
  UB1DCON_84 U38 (O[84], I[84]);
  UB1DCON_85 U39 (O[85], I[85]);
  UB1DCON_86 U40 (O[86], I[86]);
  UB1DCON_87 U41 (O[87], I[87]);
  UB1DCON_88 U42 (O[88], I[88]);
  UB1DCON_89 U43 (O[89], I[89]);
  UB1DCON_90 U44 (O[90], I[90]);
  UB1DCON_91 U45 (O[91], I[91]);
  UB1DCON_92 U46 (O[92], I[92]);
  UB1DCON_93 U47 (O[93], I[93]);
  UB1DCON_94 U48 (O[94], I[94]);
  UB1DCON_95 U49 (O[95], I[95]);
  UB1DCON_96 U50 (O[96], I[96]);
  UB1DCON_97 U51 (O[97], I[97]);
  UB1DCON_98 U52 (O[98], I[98]);
  UB1DCON_99 U53 (O[99], I[99]);
  UB1DCON_100 U54 (O[100], I[100]);
  UB1DCON_101 U55 (O[101], I[101]);
  UB1DCON_102 U56 (O[102], I[102]);
  UB1DCON_103 U57 (O[103], I[103]);
  UB1DCON_104 U58 (O[104], I[104]);
  UB1DCON_105 U59 (O[105], I[105]);
  UB1DCON_106 U60 (O[106], I[106]);
  UB1DCON_107 U61 (O[107], I[107]);
  UB1DCON_108 U62 (O[108], I[108]);
  UB1DCON_109 U63 (O[109], I[109]);
  UB1DCON_110 U64 (O[110], I[110]);
endmodule

module UBCON_111_110 (O, I);
  output [111:110] O;
  input [111:110] I;
  UB1DCON_110 U0 (O[110], I[110]);
  UB1DCON_111 U1 (O[111], I[111]);
endmodule

module UBCON_112_48 (O, I);
  output [112:48] O;
  input [112:48] I;
  UB1DCON_48 U0 (O[48], I[48]);
  UB1DCON_49 U1 (O[49], I[49]);
  UB1DCON_50 U2 (O[50], I[50]);
  UB1DCON_51 U3 (O[51], I[51]);
  UB1DCON_52 U4 (O[52], I[52]);
  UB1DCON_53 U5 (O[53], I[53]);
  UB1DCON_54 U6 (O[54], I[54]);
  UB1DCON_55 U7 (O[55], I[55]);
  UB1DCON_56 U8 (O[56], I[56]);
  UB1DCON_57 U9 (O[57], I[57]);
  UB1DCON_58 U10 (O[58], I[58]);
  UB1DCON_59 U11 (O[59], I[59]);
  UB1DCON_60 U12 (O[60], I[60]);
  UB1DCON_61 U13 (O[61], I[61]);
  UB1DCON_62 U14 (O[62], I[62]);
  UB1DCON_63 U15 (O[63], I[63]);
  UB1DCON_64 U16 (O[64], I[64]);
  UB1DCON_65 U17 (O[65], I[65]);
  UB1DCON_66 U18 (O[66], I[66]);
  UB1DCON_67 U19 (O[67], I[67]);
  UB1DCON_68 U20 (O[68], I[68]);
  UB1DCON_69 U21 (O[69], I[69]);
  UB1DCON_70 U22 (O[70], I[70]);
  UB1DCON_71 U23 (O[71], I[71]);
  UB1DCON_72 U24 (O[72], I[72]);
  UB1DCON_73 U25 (O[73], I[73]);
  UB1DCON_74 U26 (O[74], I[74]);
  UB1DCON_75 U27 (O[75], I[75]);
  UB1DCON_76 U28 (O[76], I[76]);
  UB1DCON_77 U29 (O[77], I[77]);
  UB1DCON_78 U30 (O[78], I[78]);
  UB1DCON_79 U31 (O[79], I[79]);
  UB1DCON_80 U32 (O[80], I[80]);
  UB1DCON_81 U33 (O[81], I[81]);
  UB1DCON_82 U34 (O[82], I[82]);
  UB1DCON_83 U35 (O[83], I[83]);
  UB1DCON_84 U36 (O[84], I[84]);
  UB1DCON_85 U37 (O[85], I[85]);
  UB1DCON_86 U38 (O[86], I[86]);
  UB1DCON_87 U39 (O[87], I[87]);
  UB1DCON_88 U40 (O[88], I[88]);
  UB1DCON_89 U41 (O[89], I[89]);
  UB1DCON_90 U42 (O[90], I[90]);
  UB1DCON_91 U43 (O[91], I[91]);
  UB1DCON_92 U44 (O[92], I[92]);
  UB1DCON_93 U45 (O[93], I[93]);
  UB1DCON_94 U46 (O[94], I[94]);
  UB1DCON_95 U47 (O[95], I[95]);
  UB1DCON_96 U48 (O[96], I[96]);
  UB1DCON_97 U49 (O[97], I[97]);
  UB1DCON_98 U50 (O[98], I[98]);
  UB1DCON_99 U51 (O[99], I[99]);
  UB1DCON_100 U52 (O[100], I[100]);
  UB1DCON_101 U53 (O[101], I[101]);
  UB1DCON_102 U54 (O[102], I[102]);
  UB1DCON_103 U55 (O[103], I[103]);
  UB1DCON_104 U56 (O[104], I[104]);
  UB1DCON_105 U57 (O[105], I[105]);
  UB1DCON_106 U58 (O[106], I[106]);
  UB1DCON_107 U59 (O[107], I[107]);
  UB1DCON_108 U60 (O[108], I[108]);
  UB1DCON_109 U61 (O[109], I[109]);
  UB1DCON_110 U62 (O[110], I[110]);
  UB1DCON_111 U63 (O[111], I[111]);
  UB1DCON_112 U64 (O[112], I[112]);
endmodule

module UBCON_113_112 (O, I);
  output [113:112] O;
  input [113:112] I;
  UB1DCON_112 U0 (O[112], I[112]);
  UB1DCON_113 U1 (O[113], I[113]);
endmodule

module UBCON_114_50 (O, I);
  output [114:50] O;
  input [114:50] I;
  UB1DCON_50 U0 (O[50], I[50]);
  UB1DCON_51 U1 (O[51], I[51]);
  UB1DCON_52 U2 (O[52], I[52]);
  UB1DCON_53 U3 (O[53], I[53]);
  UB1DCON_54 U4 (O[54], I[54]);
  UB1DCON_55 U5 (O[55], I[55]);
  UB1DCON_56 U6 (O[56], I[56]);
  UB1DCON_57 U7 (O[57], I[57]);
  UB1DCON_58 U8 (O[58], I[58]);
  UB1DCON_59 U9 (O[59], I[59]);
  UB1DCON_60 U10 (O[60], I[60]);
  UB1DCON_61 U11 (O[61], I[61]);
  UB1DCON_62 U12 (O[62], I[62]);
  UB1DCON_63 U13 (O[63], I[63]);
  UB1DCON_64 U14 (O[64], I[64]);
  UB1DCON_65 U15 (O[65], I[65]);
  UB1DCON_66 U16 (O[66], I[66]);
  UB1DCON_67 U17 (O[67], I[67]);
  UB1DCON_68 U18 (O[68], I[68]);
  UB1DCON_69 U19 (O[69], I[69]);
  UB1DCON_70 U20 (O[70], I[70]);
  UB1DCON_71 U21 (O[71], I[71]);
  UB1DCON_72 U22 (O[72], I[72]);
  UB1DCON_73 U23 (O[73], I[73]);
  UB1DCON_74 U24 (O[74], I[74]);
  UB1DCON_75 U25 (O[75], I[75]);
  UB1DCON_76 U26 (O[76], I[76]);
  UB1DCON_77 U27 (O[77], I[77]);
  UB1DCON_78 U28 (O[78], I[78]);
  UB1DCON_79 U29 (O[79], I[79]);
  UB1DCON_80 U30 (O[80], I[80]);
  UB1DCON_81 U31 (O[81], I[81]);
  UB1DCON_82 U32 (O[82], I[82]);
  UB1DCON_83 U33 (O[83], I[83]);
  UB1DCON_84 U34 (O[84], I[84]);
  UB1DCON_85 U35 (O[85], I[85]);
  UB1DCON_86 U36 (O[86], I[86]);
  UB1DCON_87 U37 (O[87], I[87]);
  UB1DCON_88 U38 (O[88], I[88]);
  UB1DCON_89 U39 (O[89], I[89]);
  UB1DCON_90 U40 (O[90], I[90]);
  UB1DCON_91 U41 (O[91], I[91]);
  UB1DCON_92 U42 (O[92], I[92]);
  UB1DCON_93 U43 (O[93], I[93]);
  UB1DCON_94 U44 (O[94], I[94]);
  UB1DCON_95 U45 (O[95], I[95]);
  UB1DCON_96 U46 (O[96], I[96]);
  UB1DCON_97 U47 (O[97], I[97]);
  UB1DCON_98 U48 (O[98], I[98]);
  UB1DCON_99 U49 (O[99], I[99]);
  UB1DCON_100 U50 (O[100], I[100]);
  UB1DCON_101 U51 (O[101], I[101]);
  UB1DCON_102 U52 (O[102], I[102]);
  UB1DCON_103 U53 (O[103], I[103]);
  UB1DCON_104 U54 (O[104], I[104]);
  UB1DCON_105 U55 (O[105], I[105]);
  UB1DCON_106 U56 (O[106], I[106]);
  UB1DCON_107 U57 (O[107], I[107]);
  UB1DCON_108 U58 (O[108], I[108]);
  UB1DCON_109 U59 (O[109], I[109]);
  UB1DCON_110 U60 (O[110], I[110]);
  UB1DCON_111 U61 (O[111], I[111]);
  UB1DCON_112 U62 (O[112], I[112]);
  UB1DCON_113 U63 (O[113], I[113]);
  UB1DCON_114 U64 (O[114], I[114]);
endmodule

module UBCON_115_114 (O, I);
  output [115:114] O;
  input [115:114] I;
  UB1DCON_114 U0 (O[114], I[114]);
  UB1DCON_115 U1 (O[115], I[115]);
endmodule

module UBCON_116_52 (O, I);
  output [116:52] O;
  input [116:52] I;
  UB1DCON_52 U0 (O[52], I[52]);
  UB1DCON_53 U1 (O[53], I[53]);
  UB1DCON_54 U2 (O[54], I[54]);
  UB1DCON_55 U3 (O[55], I[55]);
  UB1DCON_56 U4 (O[56], I[56]);
  UB1DCON_57 U5 (O[57], I[57]);
  UB1DCON_58 U6 (O[58], I[58]);
  UB1DCON_59 U7 (O[59], I[59]);
  UB1DCON_60 U8 (O[60], I[60]);
  UB1DCON_61 U9 (O[61], I[61]);
  UB1DCON_62 U10 (O[62], I[62]);
  UB1DCON_63 U11 (O[63], I[63]);
  UB1DCON_64 U12 (O[64], I[64]);
  UB1DCON_65 U13 (O[65], I[65]);
  UB1DCON_66 U14 (O[66], I[66]);
  UB1DCON_67 U15 (O[67], I[67]);
  UB1DCON_68 U16 (O[68], I[68]);
  UB1DCON_69 U17 (O[69], I[69]);
  UB1DCON_70 U18 (O[70], I[70]);
  UB1DCON_71 U19 (O[71], I[71]);
  UB1DCON_72 U20 (O[72], I[72]);
  UB1DCON_73 U21 (O[73], I[73]);
  UB1DCON_74 U22 (O[74], I[74]);
  UB1DCON_75 U23 (O[75], I[75]);
  UB1DCON_76 U24 (O[76], I[76]);
  UB1DCON_77 U25 (O[77], I[77]);
  UB1DCON_78 U26 (O[78], I[78]);
  UB1DCON_79 U27 (O[79], I[79]);
  UB1DCON_80 U28 (O[80], I[80]);
  UB1DCON_81 U29 (O[81], I[81]);
  UB1DCON_82 U30 (O[82], I[82]);
  UB1DCON_83 U31 (O[83], I[83]);
  UB1DCON_84 U32 (O[84], I[84]);
  UB1DCON_85 U33 (O[85], I[85]);
  UB1DCON_86 U34 (O[86], I[86]);
  UB1DCON_87 U35 (O[87], I[87]);
  UB1DCON_88 U36 (O[88], I[88]);
  UB1DCON_89 U37 (O[89], I[89]);
  UB1DCON_90 U38 (O[90], I[90]);
  UB1DCON_91 U39 (O[91], I[91]);
  UB1DCON_92 U40 (O[92], I[92]);
  UB1DCON_93 U41 (O[93], I[93]);
  UB1DCON_94 U42 (O[94], I[94]);
  UB1DCON_95 U43 (O[95], I[95]);
  UB1DCON_96 U44 (O[96], I[96]);
  UB1DCON_97 U45 (O[97], I[97]);
  UB1DCON_98 U46 (O[98], I[98]);
  UB1DCON_99 U47 (O[99], I[99]);
  UB1DCON_100 U48 (O[100], I[100]);
  UB1DCON_101 U49 (O[101], I[101]);
  UB1DCON_102 U50 (O[102], I[102]);
  UB1DCON_103 U51 (O[103], I[103]);
  UB1DCON_104 U52 (O[104], I[104]);
  UB1DCON_105 U53 (O[105], I[105]);
  UB1DCON_106 U54 (O[106], I[106]);
  UB1DCON_107 U55 (O[107], I[107]);
  UB1DCON_108 U56 (O[108], I[108]);
  UB1DCON_109 U57 (O[109], I[109]);
  UB1DCON_110 U58 (O[110], I[110]);
  UB1DCON_111 U59 (O[111], I[111]);
  UB1DCON_112 U60 (O[112], I[112]);
  UB1DCON_113 U61 (O[113], I[113]);
  UB1DCON_114 U62 (O[114], I[114]);
  UB1DCON_115 U63 (O[115], I[115]);
  UB1DCON_116 U64 (O[116], I[116]);
endmodule

module UBCON_117_116 (O, I);
  output [117:116] O;
  input [117:116] I;
  UB1DCON_116 U0 (O[116], I[116]);
  UB1DCON_117 U1 (O[117], I[117]);
endmodule

module UBCON_118_54 (O, I);
  output [118:54] O;
  input [118:54] I;
  UB1DCON_54 U0 (O[54], I[54]);
  UB1DCON_55 U1 (O[55], I[55]);
  UB1DCON_56 U2 (O[56], I[56]);
  UB1DCON_57 U3 (O[57], I[57]);
  UB1DCON_58 U4 (O[58], I[58]);
  UB1DCON_59 U5 (O[59], I[59]);
  UB1DCON_60 U6 (O[60], I[60]);
  UB1DCON_61 U7 (O[61], I[61]);
  UB1DCON_62 U8 (O[62], I[62]);
  UB1DCON_63 U9 (O[63], I[63]);
  UB1DCON_64 U10 (O[64], I[64]);
  UB1DCON_65 U11 (O[65], I[65]);
  UB1DCON_66 U12 (O[66], I[66]);
  UB1DCON_67 U13 (O[67], I[67]);
  UB1DCON_68 U14 (O[68], I[68]);
  UB1DCON_69 U15 (O[69], I[69]);
  UB1DCON_70 U16 (O[70], I[70]);
  UB1DCON_71 U17 (O[71], I[71]);
  UB1DCON_72 U18 (O[72], I[72]);
  UB1DCON_73 U19 (O[73], I[73]);
  UB1DCON_74 U20 (O[74], I[74]);
  UB1DCON_75 U21 (O[75], I[75]);
  UB1DCON_76 U22 (O[76], I[76]);
  UB1DCON_77 U23 (O[77], I[77]);
  UB1DCON_78 U24 (O[78], I[78]);
  UB1DCON_79 U25 (O[79], I[79]);
  UB1DCON_80 U26 (O[80], I[80]);
  UB1DCON_81 U27 (O[81], I[81]);
  UB1DCON_82 U28 (O[82], I[82]);
  UB1DCON_83 U29 (O[83], I[83]);
  UB1DCON_84 U30 (O[84], I[84]);
  UB1DCON_85 U31 (O[85], I[85]);
  UB1DCON_86 U32 (O[86], I[86]);
  UB1DCON_87 U33 (O[87], I[87]);
  UB1DCON_88 U34 (O[88], I[88]);
  UB1DCON_89 U35 (O[89], I[89]);
  UB1DCON_90 U36 (O[90], I[90]);
  UB1DCON_91 U37 (O[91], I[91]);
  UB1DCON_92 U38 (O[92], I[92]);
  UB1DCON_93 U39 (O[93], I[93]);
  UB1DCON_94 U40 (O[94], I[94]);
  UB1DCON_95 U41 (O[95], I[95]);
  UB1DCON_96 U42 (O[96], I[96]);
  UB1DCON_97 U43 (O[97], I[97]);
  UB1DCON_98 U44 (O[98], I[98]);
  UB1DCON_99 U45 (O[99], I[99]);
  UB1DCON_100 U46 (O[100], I[100]);
  UB1DCON_101 U47 (O[101], I[101]);
  UB1DCON_102 U48 (O[102], I[102]);
  UB1DCON_103 U49 (O[103], I[103]);
  UB1DCON_104 U50 (O[104], I[104]);
  UB1DCON_105 U51 (O[105], I[105]);
  UB1DCON_106 U52 (O[106], I[106]);
  UB1DCON_107 U53 (O[107], I[107]);
  UB1DCON_108 U54 (O[108], I[108]);
  UB1DCON_109 U55 (O[109], I[109]);
  UB1DCON_110 U56 (O[110], I[110]);
  UB1DCON_111 U57 (O[111], I[111]);
  UB1DCON_112 U58 (O[112], I[112]);
  UB1DCON_113 U59 (O[113], I[113]);
  UB1DCON_114 U60 (O[114], I[114]);
  UB1DCON_115 U61 (O[115], I[115]);
  UB1DCON_116 U62 (O[116], I[116]);
  UB1DCON_117 U63 (O[117], I[117]);
  UB1DCON_118 U64 (O[118], I[118]);
endmodule

module UBCON_119_116 (O, I);
  output [119:116] O;
  input [119:116] I;
  UB1DCON_116 U0 (O[116], I[116]);
  UB1DCON_117 U1 (O[117], I[117]);
  UB1DCON_118 U2 (O[118], I[118]);
  UB1DCON_119 U3 (O[119], I[119]);
endmodule

module UBCON_119_118 (O, I);
  output [119:118] O;
  input [119:118] I;
  UB1DCON_118 U0 (O[118], I[118]);
  UB1DCON_119 U1 (O[119], I[119]);
endmodule

module UBCON_11_0 (O, I);
  output [11:0] O;
  input [11:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
endmodule

module UBCON_11_10 (O, I);
  output [11:10] O;
  input [11:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
endmodule

module UBCON_11_2 (O, I);
  output [11:2] O;
  input [11:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
  UB1DCON_9 U7 (O[9], I[9]);
  UB1DCON_10 U8 (O[10], I[10]);
  UB1DCON_11 U9 (O[11], I[11]);
endmodule

module UBCON_11_4 (O, I);
  output [11:4] O;
  input [11:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
endmodule

module UBCON_11_6 (O, I);
  output [11:6] O;
  input [11:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
  UB1DCON_9 U3 (O[9], I[9]);
  UB1DCON_10 U4 (O[10], I[10]);
  UB1DCON_11 U5 (O[11], I[11]);
endmodule

module UBCON_11_8 (O, I);
  output [11:8] O;
  input [11:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
  UB1DCON_11 U3 (O[11], I[11]);
endmodule

module UBCON_120_56 (O, I);
  output [120:56] O;
  input [120:56] I;
  UB1DCON_56 U0 (O[56], I[56]);
  UB1DCON_57 U1 (O[57], I[57]);
  UB1DCON_58 U2 (O[58], I[58]);
  UB1DCON_59 U3 (O[59], I[59]);
  UB1DCON_60 U4 (O[60], I[60]);
  UB1DCON_61 U5 (O[61], I[61]);
  UB1DCON_62 U6 (O[62], I[62]);
  UB1DCON_63 U7 (O[63], I[63]);
  UB1DCON_64 U8 (O[64], I[64]);
  UB1DCON_65 U9 (O[65], I[65]);
  UB1DCON_66 U10 (O[66], I[66]);
  UB1DCON_67 U11 (O[67], I[67]);
  UB1DCON_68 U12 (O[68], I[68]);
  UB1DCON_69 U13 (O[69], I[69]);
  UB1DCON_70 U14 (O[70], I[70]);
  UB1DCON_71 U15 (O[71], I[71]);
  UB1DCON_72 U16 (O[72], I[72]);
  UB1DCON_73 U17 (O[73], I[73]);
  UB1DCON_74 U18 (O[74], I[74]);
  UB1DCON_75 U19 (O[75], I[75]);
  UB1DCON_76 U20 (O[76], I[76]);
  UB1DCON_77 U21 (O[77], I[77]);
  UB1DCON_78 U22 (O[78], I[78]);
  UB1DCON_79 U23 (O[79], I[79]);
  UB1DCON_80 U24 (O[80], I[80]);
  UB1DCON_81 U25 (O[81], I[81]);
  UB1DCON_82 U26 (O[82], I[82]);
  UB1DCON_83 U27 (O[83], I[83]);
  UB1DCON_84 U28 (O[84], I[84]);
  UB1DCON_85 U29 (O[85], I[85]);
  UB1DCON_86 U30 (O[86], I[86]);
  UB1DCON_87 U31 (O[87], I[87]);
  UB1DCON_88 U32 (O[88], I[88]);
  UB1DCON_89 U33 (O[89], I[89]);
  UB1DCON_90 U34 (O[90], I[90]);
  UB1DCON_91 U35 (O[91], I[91]);
  UB1DCON_92 U36 (O[92], I[92]);
  UB1DCON_93 U37 (O[93], I[93]);
  UB1DCON_94 U38 (O[94], I[94]);
  UB1DCON_95 U39 (O[95], I[95]);
  UB1DCON_96 U40 (O[96], I[96]);
  UB1DCON_97 U41 (O[97], I[97]);
  UB1DCON_98 U42 (O[98], I[98]);
  UB1DCON_99 U43 (O[99], I[99]);
  UB1DCON_100 U44 (O[100], I[100]);
  UB1DCON_101 U45 (O[101], I[101]);
  UB1DCON_102 U46 (O[102], I[102]);
  UB1DCON_103 U47 (O[103], I[103]);
  UB1DCON_104 U48 (O[104], I[104]);
  UB1DCON_105 U49 (O[105], I[105]);
  UB1DCON_106 U50 (O[106], I[106]);
  UB1DCON_107 U51 (O[107], I[107]);
  UB1DCON_108 U52 (O[108], I[108]);
  UB1DCON_109 U53 (O[109], I[109]);
  UB1DCON_110 U54 (O[110], I[110]);
  UB1DCON_111 U55 (O[111], I[111]);
  UB1DCON_112 U56 (O[112], I[112]);
  UB1DCON_113 U57 (O[113], I[113]);
  UB1DCON_114 U58 (O[114], I[114]);
  UB1DCON_115 U59 (O[115], I[115]);
  UB1DCON_116 U60 (O[116], I[116]);
  UB1DCON_117 U61 (O[117], I[117]);
  UB1DCON_118 U62 (O[118], I[118]);
  UB1DCON_119 U63 (O[119], I[119]);
  UB1DCON_120 U64 (O[120], I[120]);
endmodule

module UBCON_121_116 (O, I);
  output [121:116] O;
  input [121:116] I;
  UB1DCON_116 U0 (O[116], I[116]);
  UB1DCON_117 U1 (O[117], I[117]);
  UB1DCON_118 U2 (O[118], I[118]);
  UB1DCON_119 U3 (O[119], I[119]);
  UB1DCON_120 U4 (O[120], I[120]);
  UB1DCON_121 U5 (O[121], I[121]);
endmodule

module UBCON_121_120 (O, I);
  output [121:120] O;
  input [121:120] I;
  UB1DCON_120 U0 (O[120], I[120]);
  UB1DCON_121 U1 (O[121], I[121]);
endmodule

module UBCON_122_58 (O, I);
  output [122:58] O;
  input [122:58] I;
  UB1DCON_58 U0 (O[58], I[58]);
  UB1DCON_59 U1 (O[59], I[59]);
  UB1DCON_60 U2 (O[60], I[60]);
  UB1DCON_61 U3 (O[61], I[61]);
  UB1DCON_62 U4 (O[62], I[62]);
  UB1DCON_63 U5 (O[63], I[63]);
  UB1DCON_64 U6 (O[64], I[64]);
  UB1DCON_65 U7 (O[65], I[65]);
  UB1DCON_66 U8 (O[66], I[66]);
  UB1DCON_67 U9 (O[67], I[67]);
  UB1DCON_68 U10 (O[68], I[68]);
  UB1DCON_69 U11 (O[69], I[69]);
  UB1DCON_70 U12 (O[70], I[70]);
  UB1DCON_71 U13 (O[71], I[71]);
  UB1DCON_72 U14 (O[72], I[72]);
  UB1DCON_73 U15 (O[73], I[73]);
  UB1DCON_74 U16 (O[74], I[74]);
  UB1DCON_75 U17 (O[75], I[75]);
  UB1DCON_76 U18 (O[76], I[76]);
  UB1DCON_77 U19 (O[77], I[77]);
  UB1DCON_78 U20 (O[78], I[78]);
  UB1DCON_79 U21 (O[79], I[79]);
  UB1DCON_80 U22 (O[80], I[80]);
  UB1DCON_81 U23 (O[81], I[81]);
  UB1DCON_82 U24 (O[82], I[82]);
  UB1DCON_83 U25 (O[83], I[83]);
  UB1DCON_84 U26 (O[84], I[84]);
  UB1DCON_85 U27 (O[85], I[85]);
  UB1DCON_86 U28 (O[86], I[86]);
  UB1DCON_87 U29 (O[87], I[87]);
  UB1DCON_88 U30 (O[88], I[88]);
  UB1DCON_89 U31 (O[89], I[89]);
  UB1DCON_90 U32 (O[90], I[90]);
  UB1DCON_91 U33 (O[91], I[91]);
  UB1DCON_92 U34 (O[92], I[92]);
  UB1DCON_93 U35 (O[93], I[93]);
  UB1DCON_94 U36 (O[94], I[94]);
  UB1DCON_95 U37 (O[95], I[95]);
  UB1DCON_96 U38 (O[96], I[96]);
  UB1DCON_97 U39 (O[97], I[97]);
  UB1DCON_98 U40 (O[98], I[98]);
  UB1DCON_99 U41 (O[99], I[99]);
  UB1DCON_100 U42 (O[100], I[100]);
  UB1DCON_101 U43 (O[101], I[101]);
  UB1DCON_102 U44 (O[102], I[102]);
  UB1DCON_103 U45 (O[103], I[103]);
  UB1DCON_104 U46 (O[104], I[104]);
  UB1DCON_105 U47 (O[105], I[105]);
  UB1DCON_106 U48 (O[106], I[106]);
  UB1DCON_107 U49 (O[107], I[107]);
  UB1DCON_108 U50 (O[108], I[108]);
  UB1DCON_109 U51 (O[109], I[109]);
  UB1DCON_110 U52 (O[110], I[110]);
  UB1DCON_111 U53 (O[111], I[111]);
  UB1DCON_112 U54 (O[112], I[112]);
  UB1DCON_113 U55 (O[113], I[113]);
  UB1DCON_114 U56 (O[114], I[114]);
  UB1DCON_115 U57 (O[115], I[115]);
  UB1DCON_116 U58 (O[116], I[116]);
  UB1DCON_117 U59 (O[117], I[117]);
  UB1DCON_118 U60 (O[118], I[118]);
  UB1DCON_119 U61 (O[119], I[119]);
  UB1DCON_120 U62 (O[120], I[120]);
  UB1DCON_121 U63 (O[121], I[121]);
  UB1DCON_122 U64 (O[122], I[122]);
endmodule

module UBCON_123_116 (O, I);
  output [123:116] O;
  input [123:116] I;
  UB1DCON_116 U0 (O[116], I[116]);
  UB1DCON_117 U1 (O[117], I[117]);
  UB1DCON_118 U2 (O[118], I[118]);
  UB1DCON_119 U3 (O[119], I[119]);
  UB1DCON_120 U4 (O[120], I[120]);
  UB1DCON_121 U5 (O[121], I[121]);
  UB1DCON_122 U6 (O[122], I[122]);
  UB1DCON_123 U7 (O[123], I[123]);
endmodule

module UBCON_123_122 (O, I);
  output [123:122] O;
  input [123:122] I;
  UB1DCON_122 U0 (O[122], I[122]);
  UB1DCON_123 U1 (O[123], I[123]);
endmodule

module UBCON_124_60 (O, I);
  output [124:60] O;
  input [124:60] I;
  UB1DCON_60 U0 (O[60], I[60]);
  UB1DCON_61 U1 (O[61], I[61]);
  UB1DCON_62 U2 (O[62], I[62]);
  UB1DCON_63 U3 (O[63], I[63]);
  UB1DCON_64 U4 (O[64], I[64]);
  UB1DCON_65 U5 (O[65], I[65]);
  UB1DCON_66 U6 (O[66], I[66]);
  UB1DCON_67 U7 (O[67], I[67]);
  UB1DCON_68 U8 (O[68], I[68]);
  UB1DCON_69 U9 (O[69], I[69]);
  UB1DCON_70 U10 (O[70], I[70]);
  UB1DCON_71 U11 (O[71], I[71]);
  UB1DCON_72 U12 (O[72], I[72]);
  UB1DCON_73 U13 (O[73], I[73]);
  UB1DCON_74 U14 (O[74], I[74]);
  UB1DCON_75 U15 (O[75], I[75]);
  UB1DCON_76 U16 (O[76], I[76]);
  UB1DCON_77 U17 (O[77], I[77]);
  UB1DCON_78 U18 (O[78], I[78]);
  UB1DCON_79 U19 (O[79], I[79]);
  UB1DCON_80 U20 (O[80], I[80]);
  UB1DCON_81 U21 (O[81], I[81]);
  UB1DCON_82 U22 (O[82], I[82]);
  UB1DCON_83 U23 (O[83], I[83]);
  UB1DCON_84 U24 (O[84], I[84]);
  UB1DCON_85 U25 (O[85], I[85]);
  UB1DCON_86 U26 (O[86], I[86]);
  UB1DCON_87 U27 (O[87], I[87]);
  UB1DCON_88 U28 (O[88], I[88]);
  UB1DCON_89 U29 (O[89], I[89]);
  UB1DCON_90 U30 (O[90], I[90]);
  UB1DCON_91 U31 (O[91], I[91]);
  UB1DCON_92 U32 (O[92], I[92]);
  UB1DCON_93 U33 (O[93], I[93]);
  UB1DCON_94 U34 (O[94], I[94]);
  UB1DCON_95 U35 (O[95], I[95]);
  UB1DCON_96 U36 (O[96], I[96]);
  UB1DCON_97 U37 (O[97], I[97]);
  UB1DCON_98 U38 (O[98], I[98]);
  UB1DCON_99 U39 (O[99], I[99]);
  UB1DCON_100 U40 (O[100], I[100]);
  UB1DCON_101 U41 (O[101], I[101]);
  UB1DCON_102 U42 (O[102], I[102]);
  UB1DCON_103 U43 (O[103], I[103]);
  UB1DCON_104 U44 (O[104], I[104]);
  UB1DCON_105 U45 (O[105], I[105]);
  UB1DCON_106 U46 (O[106], I[106]);
  UB1DCON_107 U47 (O[107], I[107]);
  UB1DCON_108 U48 (O[108], I[108]);
  UB1DCON_109 U49 (O[109], I[109]);
  UB1DCON_110 U50 (O[110], I[110]);
  UB1DCON_111 U51 (O[111], I[111]);
  UB1DCON_112 U52 (O[112], I[112]);
  UB1DCON_113 U53 (O[113], I[113]);
  UB1DCON_114 U54 (O[114], I[114]);
  UB1DCON_115 U55 (O[115], I[115]);
  UB1DCON_116 U56 (O[116], I[116]);
  UB1DCON_117 U57 (O[117], I[117]);
  UB1DCON_118 U58 (O[118], I[118]);
  UB1DCON_119 U59 (O[119], I[119]);
  UB1DCON_120 U60 (O[120], I[120]);
  UB1DCON_121 U61 (O[121], I[121]);
  UB1DCON_122 U62 (O[122], I[122]);
  UB1DCON_123 U63 (O[123], I[123]);
  UB1DCON_124 U64 (O[124], I[124]);
endmodule

module UBCON_125_116 (O, I);
  output [125:116] O;
  input [125:116] I;
  UB1DCON_116 U0 (O[116], I[116]);
  UB1DCON_117 U1 (O[117], I[117]);
  UB1DCON_118 U2 (O[118], I[118]);
  UB1DCON_119 U3 (O[119], I[119]);
  UB1DCON_120 U4 (O[120], I[120]);
  UB1DCON_121 U5 (O[121], I[121]);
  UB1DCON_122 U6 (O[122], I[122]);
  UB1DCON_123 U7 (O[123], I[123]);
  UB1DCON_124 U8 (O[124], I[124]);
  UB1DCON_125 U9 (O[125], I[125]);
endmodule

module UBCON_125_124 (O, I);
  output [125:124] O;
  input [125:124] I;
  UB1DCON_124 U0 (O[124], I[124]);
  UB1DCON_125 U1 (O[125], I[125]);
endmodule

module UBCON_126_0 (O, I);
  output [126:0] O;
  input [126:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
  UB1DCON_28 U28 (O[28], I[28]);
  UB1DCON_29 U29 (O[29], I[29]);
  UB1DCON_30 U30 (O[30], I[30]);
  UB1DCON_31 U31 (O[31], I[31]);
  UB1DCON_32 U32 (O[32], I[32]);
  UB1DCON_33 U33 (O[33], I[33]);
  UB1DCON_34 U34 (O[34], I[34]);
  UB1DCON_35 U35 (O[35], I[35]);
  UB1DCON_36 U36 (O[36], I[36]);
  UB1DCON_37 U37 (O[37], I[37]);
  UB1DCON_38 U38 (O[38], I[38]);
  UB1DCON_39 U39 (O[39], I[39]);
  UB1DCON_40 U40 (O[40], I[40]);
  UB1DCON_41 U41 (O[41], I[41]);
  UB1DCON_42 U42 (O[42], I[42]);
  UB1DCON_43 U43 (O[43], I[43]);
  UB1DCON_44 U44 (O[44], I[44]);
  UB1DCON_45 U45 (O[45], I[45]);
  UB1DCON_46 U46 (O[46], I[46]);
  UB1DCON_47 U47 (O[47], I[47]);
  UB1DCON_48 U48 (O[48], I[48]);
  UB1DCON_49 U49 (O[49], I[49]);
  UB1DCON_50 U50 (O[50], I[50]);
  UB1DCON_51 U51 (O[51], I[51]);
  UB1DCON_52 U52 (O[52], I[52]);
  UB1DCON_53 U53 (O[53], I[53]);
  UB1DCON_54 U54 (O[54], I[54]);
  UB1DCON_55 U55 (O[55], I[55]);
  UB1DCON_56 U56 (O[56], I[56]);
  UB1DCON_57 U57 (O[57], I[57]);
  UB1DCON_58 U58 (O[58], I[58]);
  UB1DCON_59 U59 (O[59], I[59]);
  UB1DCON_60 U60 (O[60], I[60]);
  UB1DCON_61 U61 (O[61], I[61]);
  UB1DCON_62 U62 (O[62], I[62]);
  UB1DCON_63 U63 (O[63], I[63]);
  UB1DCON_64 U64 (O[64], I[64]);
  UB1DCON_65 U65 (O[65], I[65]);
  UB1DCON_66 U66 (O[66], I[66]);
  UB1DCON_67 U67 (O[67], I[67]);
  UB1DCON_68 U68 (O[68], I[68]);
  UB1DCON_69 U69 (O[69], I[69]);
  UB1DCON_70 U70 (O[70], I[70]);
  UB1DCON_71 U71 (O[71], I[71]);
  UB1DCON_72 U72 (O[72], I[72]);
  UB1DCON_73 U73 (O[73], I[73]);
  UB1DCON_74 U74 (O[74], I[74]);
  UB1DCON_75 U75 (O[75], I[75]);
  UB1DCON_76 U76 (O[76], I[76]);
  UB1DCON_77 U77 (O[77], I[77]);
  UB1DCON_78 U78 (O[78], I[78]);
  UB1DCON_79 U79 (O[79], I[79]);
  UB1DCON_80 U80 (O[80], I[80]);
  UB1DCON_81 U81 (O[81], I[81]);
  UB1DCON_82 U82 (O[82], I[82]);
  UB1DCON_83 U83 (O[83], I[83]);
  UB1DCON_84 U84 (O[84], I[84]);
  UB1DCON_85 U85 (O[85], I[85]);
  UB1DCON_86 U86 (O[86], I[86]);
  UB1DCON_87 U87 (O[87], I[87]);
  UB1DCON_88 U88 (O[88], I[88]);
  UB1DCON_89 U89 (O[89], I[89]);
  UB1DCON_90 U90 (O[90], I[90]);
  UB1DCON_91 U91 (O[91], I[91]);
  UB1DCON_92 U92 (O[92], I[92]);
  UB1DCON_93 U93 (O[93], I[93]);
  UB1DCON_94 U94 (O[94], I[94]);
  UB1DCON_95 U95 (O[95], I[95]);
  UB1DCON_96 U96 (O[96], I[96]);
  UB1DCON_97 U97 (O[97], I[97]);
  UB1DCON_98 U98 (O[98], I[98]);
  UB1DCON_99 U99 (O[99], I[99]);
  UB1DCON_100 U100 (O[100], I[100]);
  UB1DCON_101 U101 (O[101], I[101]);
  UB1DCON_102 U102 (O[102], I[102]);
  UB1DCON_103 U103 (O[103], I[103]);
  UB1DCON_104 U104 (O[104], I[104]);
  UB1DCON_105 U105 (O[105], I[105]);
  UB1DCON_106 U106 (O[106], I[106]);
  UB1DCON_107 U107 (O[107], I[107]);
  UB1DCON_108 U108 (O[108], I[108]);
  UB1DCON_109 U109 (O[109], I[109]);
  UB1DCON_110 U110 (O[110], I[110]);
  UB1DCON_111 U111 (O[111], I[111]);
  UB1DCON_112 U112 (O[112], I[112]);
  UB1DCON_113 U113 (O[113], I[113]);
  UB1DCON_114 U114 (O[114], I[114]);
  UB1DCON_115 U115 (O[115], I[115]);
  UB1DCON_116 U116 (O[116], I[116]);
  UB1DCON_117 U117 (O[117], I[117]);
  UB1DCON_118 U118 (O[118], I[118]);
  UB1DCON_119 U119 (O[119], I[119]);
  UB1DCON_120 U120 (O[120], I[120]);
  UB1DCON_121 U121 (O[121], I[121]);
  UB1DCON_122 U122 (O[122], I[122]);
  UB1DCON_123 U123 (O[123], I[123]);
  UB1DCON_124 U124 (O[124], I[124]);
  UB1DCON_125 U125 (O[125], I[125]);
  UB1DCON_126 U126 (O[126], I[126]);
endmodule

module UBCON_126_116 (O, I);
  output [126:116] O;
  input [126:116] I;
  UB1DCON_116 U0 (O[116], I[116]);
  UB1DCON_117 U1 (O[117], I[117]);
  UB1DCON_118 U2 (O[118], I[118]);
  UB1DCON_119 U3 (O[119], I[119]);
  UB1DCON_120 U4 (O[120], I[120]);
  UB1DCON_121 U5 (O[121], I[121]);
  UB1DCON_122 U6 (O[122], I[122]);
  UB1DCON_123 U7 (O[123], I[123]);
  UB1DCON_124 U8 (O[124], I[124]);
  UB1DCON_125 U9 (O[125], I[125]);
  UB1DCON_126 U10 (O[126], I[126]);
endmodule

module UBCON_126_124 (O, I);
  output [126:124] O;
  input [126:124] I;
  UB1DCON_124 U0 (O[124], I[124]);
  UB1DCON_125 U1 (O[125], I[125]);
  UB1DCON_126 U2 (O[126], I[126]);
endmodule

module UBCON_126_62 (O, I);
  output [126:62] O;
  input [126:62] I;
  UB1DCON_62 U0 (O[62], I[62]);
  UB1DCON_63 U1 (O[63], I[63]);
  UB1DCON_64 U2 (O[64], I[64]);
  UB1DCON_65 U3 (O[65], I[65]);
  UB1DCON_66 U4 (O[66], I[66]);
  UB1DCON_67 U5 (O[67], I[67]);
  UB1DCON_68 U6 (O[68], I[68]);
  UB1DCON_69 U7 (O[69], I[69]);
  UB1DCON_70 U8 (O[70], I[70]);
  UB1DCON_71 U9 (O[71], I[71]);
  UB1DCON_72 U10 (O[72], I[72]);
  UB1DCON_73 U11 (O[73], I[73]);
  UB1DCON_74 U12 (O[74], I[74]);
  UB1DCON_75 U13 (O[75], I[75]);
  UB1DCON_76 U14 (O[76], I[76]);
  UB1DCON_77 U15 (O[77], I[77]);
  UB1DCON_78 U16 (O[78], I[78]);
  UB1DCON_79 U17 (O[79], I[79]);
  UB1DCON_80 U18 (O[80], I[80]);
  UB1DCON_81 U19 (O[81], I[81]);
  UB1DCON_82 U20 (O[82], I[82]);
  UB1DCON_83 U21 (O[83], I[83]);
  UB1DCON_84 U22 (O[84], I[84]);
  UB1DCON_85 U23 (O[85], I[85]);
  UB1DCON_86 U24 (O[86], I[86]);
  UB1DCON_87 U25 (O[87], I[87]);
  UB1DCON_88 U26 (O[88], I[88]);
  UB1DCON_89 U27 (O[89], I[89]);
  UB1DCON_90 U28 (O[90], I[90]);
  UB1DCON_91 U29 (O[91], I[91]);
  UB1DCON_92 U30 (O[92], I[92]);
  UB1DCON_93 U31 (O[93], I[93]);
  UB1DCON_94 U32 (O[94], I[94]);
  UB1DCON_95 U33 (O[95], I[95]);
  UB1DCON_96 U34 (O[96], I[96]);
  UB1DCON_97 U35 (O[97], I[97]);
  UB1DCON_98 U36 (O[98], I[98]);
  UB1DCON_99 U37 (O[99], I[99]);
  UB1DCON_100 U38 (O[100], I[100]);
  UB1DCON_101 U39 (O[101], I[101]);
  UB1DCON_102 U40 (O[102], I[102]);
  UB1DCON_103 U41 (O[103], I[103]);
  UB1DCON_104 U42 (O[104], I[104]);
  UB1DCON_105 U43 (O[105], I[105]);
  UB1DCON_106 U44 (O[106], I[106]);
  UB1DCON_107 U45 (O[107], I[107]);
  UB1DCON_108 U46 (O[108], I[108]);
  UB1DCON_109 U47 (O[109], I[109]);
  UB1DCON_110 U48 (O[110], I[110]);
  UB1DCON_111 U49 (O[111], I[111]);
  UB1DCON_112 U50 (O[112], I[112]);
  UB1DCON_113 U51 (O[113], I[113]);
  UB1DCON_114 U52 (O[114], I[114]);
  UB1DCON_115 U53 (O[115], I[115]);
  UB1DCON_116 U54 (O[116], I[116]);
  UB1DCON_117 U55 (O[117], I[117]);
  UB1DCON_118 U56 (O[118], I[118]);
  UB1DCON_119 U57 (O[119], I[119]);
  UB1DCON_120 U58 (O[120], I[120]);
  UB1DCON_121 U59 (O[121], I[121]);
  UB1DCON_122 U60 (O[122], I[122]);
  UB1DCON_123 U61 (O[123], I[123]);
  UB1DCON_124 U62 (O[124], I[124]);
  UB1DCON_125 U63 (O[125], I[125]);
  UB1DCON_126 U64 (O[126], I[126]);
endmodule

module UBCON_15_14 (O, I);
  output [15:14] O;
  input [15:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
endmodule

module UBCON_17_16 (O, I);
  output [17:16] O;
  input [17:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
endmodule

module UBCON_19_18 (O, I);
  output [19:18] O;
  input [19:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_23_22 (O, I);
  output [23:22] O;
  input [23:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
endmodule

module UBCON_25_24 (O, I);
  output [25:24] O;
  input [25:24] I;
  UB1DCON_24 U0 (O[24], I[24]);
  UB1DCON_25 U1 (O[25], I[25]);
endmodule

module UBCON_27_0 (O, I);
  output [27:0] O;
  input [27:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
endmodule

module UBCON_27_10 (O, I);
  output [27:10] O;
  input [27:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
  UB1DCON_13 U3 (O[13], I[13]);
  UB1DCON_14 U4 (O[14], I[14]);
  UB1DCON_15 U5 (O[15], I[15]);
  UB1DCON_16 U6 (O[16], I[16]);
  UB1DCON_17 U7 (O[17], I[17]);
  UB1DCON_18 U8 (O[18], I[18]);
  UB1DCON_19 U9 (O[19], I[19]);
  UB1DCON_20 U10 (O[20], I[20]);
  UB1DCON_21 U11 (O[21], I[21]);
  UB1DCON_22 U12 (O[22], I[22]);
  UB1DCON_23 U13 (O[23], I[23]);
  UB1DCON_24 U14 (O[24], I[24]);
  UB1DCON_25 U15 (O[25], I[25]);
  UB1DCON_26 U16 (O[26], I[26]);
  UB1DCON_27 U17 (O[27], I[27]);
endmodule

module UBCON_27_12 (O, I);
  output [27:12] O;
  input [27:12] I;
  UB1DCON_12 U0 (O[12], I[12]);
  UB1DCON_13 U1 (O[13], I[13]);
  UB1DCON_14 U2 (O[14], I[14]);
  UB1DCON_15 U3 (O[15], I[15]);
  UB1DCON_16 U4 (O[16], I[16]);
  UB1DCON_17 U5 (O[17], I[17]);
  UB1DCON_18 U6 (O[18], I[18]);
  UB1DCON_19 U7 (O[19], I[19]);
  UB1DCON_20 U8 (O[20], I[20]);
  UB1DCON_21 U9 (O[21], I[21]);
  UB1DCON_22 U10 (O[22], I[22]);
  UB1DCON_23 U11 (O[23], I[23]);
  UB1DCON_24 U12 (O[24], I[24]);
  UB1DCON_25 U13 (O[25], I[25]);
  UB1DCON_26 U14 (O[26], I[26]);
  UB1DCON_27 U15 (O[27], I[27]);
endmodule

module UBCON_27_14 (O, I);
  output [27:14] O;
  input [27:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
  UB1DCON_18 U4 (O[18], I[18]);
  UB1DCON_19 U5 (O[19], I[19]);
  UB1DCON_20 U6 (O[20], I[20]);
  UB1DCON_21 U7 (O[21], I[21]);
  UB1DCON_22 U8 (O[22], I[22]);
  UB1DCON_23 U9 (O[23], I[23]);
  UB1DCON_24 U10 (O[24], I[24]);
  UB1DCON_25 U11 (O[25], I[25]);
  UB1DCON_26 U12 (O[26], I[26]);
  UB1DCON_27 U13 (O[27], I[27]);
endmodule

module UBCON_27_16 (O, I);
  output [27:16] O;
  input [27:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
  UB1DCON_19 U3 (O[19], I[19]);
  UB1DCON_20 U4 (O[20], I[20]);
  UB1DCON_21 U5 (O[21], I[21]);
  UB1DCON_22 U6 (O[22], I[22]);
  UB1DCON_23 U7 (O[23], I[23]);
  UB1DCON_24 U8 (O[24], I[24]);
  UB1DCON_25 U9 (O[25], I[25]);
  UB1DCON_26 U10 (O[26], I[26]);
  UB1DCON_27 U11 (O[27], I[27]);
endmodule

module UBCON_27_18 (O, I);
  output [27:18] O;
  input [27:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
  UB1DCON_20 U2 (O[20], I[20]);
  UB1DCON_21 U3 (O[21], I[21]);
  UB1DCON_22 U4 (O[22], I[22]);
  UB1DCON_23 U5 (O[23], I[23]);
  UB1DCON_24 U6 (O[24], I[24]);
  UB1DCON_25 U7 (O[25], I[25]);
  UB1DCON_26 U8 (O[26], I[26]);
  UB1DCON_27 U9 (O[27], I[27]);
endmodule

module UBCON_27_2 (O, I);
  output [27:2] O;
  input [27:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
  UB1DCON_9 U7 (O[9], I[9]);
  UB1DCON_10 U8 (O[10], I[10]);
  UB1DCON_11 U9 (O[11], I[11]);
  UB1DCON_12 U10 (O[12], I[12]);
  UB1DCON_13 U11 (O[13], I[13]);
  UB1DCON_14 U12 (O[14], I[14]);
  UB1DCON_15 U13 (O[15], I[15]);
  UB1DCON_16 U14 (O[16], I[16]);
  UB1DCON_17 U15 (O[17], I[17]);
  UB1DCON_18 U16 (O[18], I[18]);
  UB1DCON_19 U17 (O[19], I[19]);
  UB1DCON_20 U18 (O[20], I[20]);
  UB1DCON_21 U19 (O[21], I[21]);
  UB1DCON_22 U20 (O[22], I[22]);
  UB1DCON_23 U21 (O[23], I[23]);
  UB1DCON_24 U22 (O[24], I[24]);
  UB1DCON_25 U23 (O[25], I[25]);
  UB1DCON_26 U24 (O[26], I[26]);
  UB1DCON_27 U25 (O[27], I[27]);
endmodule

module UBCON_27_20 (O, I);
  output [27:20] O;
  input [27:20] I;
  UB1DCON_20 U0 (O[20], I[20]);
  UB1DCON_21 U1 (O[21], I[21]);
  UB1DCON_22 U2 (O[22], I[22]);
  UB1DCON_23 U3 (O[23], I[23]);
  UB1DCON_24 U4 (O[24], I[24]);
  UB1DCON_25 U5 (O[25], I[25]);
  UB1DCON_26 U6 (O[26], I[26]);
  UB1DCON_27 U7 (O[27], I[27]);
endmodule

module UBCON_27_22 (O, I);
  output [27:22] O;
  input [27:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
  UB1DCON_24 U2 (O[24], I[24]);
  UB1DCON_25 U3 (O[25], I[25]);
  UB1DCON_26 U4 (O[26], I[26]);
  UB1DCON_27 U5 (O[27], I[27]);
endmodule

module UBCON_27_24 (O, I);
  output [27:24] O;
  input [27:24] I;
  UB1DCON_24 U0 (O[24], I[24]);
  UB1DCON_25 U1 (O[25], I[25]);
  UB1DCON_26 U2 (O[26], I[26]);
  UB1DCON_27 U3 (O[27], I[27]);
endmodule

module UBCON_27_26 (O, I);
  output [27:26] O;
  input [27:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
endmodule

module UBCON_27_4 (O, I);
  output [27:4] O;
  input [27:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
  UB1DCON_19 U15 (O[19], I[19]);
  UB1DCON_20 U16 (O[20], I[20]);
  UB1DCON_21 U17 (O[21], I[21]);
  UB1DCON_22 U18 (O[22], I[22]);
  UB1DCON_23 U19 (O[23], I[23]);
  UB1DCON_24 U20 (O[24], I[24]);
  UB1DCON_25 U21 (O[25], I[25]);
  UB1DCON_26 U22 (O[26], I[26]);
  UB1DCON_27 U23 (O[27], I[27]);
endmodule

module UBCON_27_6 (O, I);
  output [27:6] O;
  input [27:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
  UB1DCON_9 U3 (O[9], I[9]);
  UB1DCON_10 U4 (O[10], I[10]);
  UB1DCON_11 U5 (O[11], I[11]);
  UB1DCON_12 U6 (O[12], I[12]);
  UB1DCON_13 U7 (O[13], I[13]);
  UB1DCON_14 U8 (O[14], I[14]);
  UB1DCON_15 U9 (O[15], I[15]);
  UB1DCON_16 U10 (O[16], I[16]);
  UB1DCON_17 U11 (O[17], I[17]);
  UB1DCON_18 U12 (O[18], I[18]);
  UB1DCON_19 U13 (O[19], I[19]);
  UB1DCON_20 U14 (O[20], I[20]);
  UB1DCON_21 U15 (O[21], I[21]);
  UB1DCON_22 U16 (O[22], I[22]);
  UB1DCON_23 U17 (O[23], I[23]);
  UB1DCON_24 U18 (O[24], I[24]);
  UB1DCON_25 U19 (O[25], I[25]);
  UB1DCON_26 U20 (O[26], I[26]);
  UB1DCON_27 U21 (O[27], I[27]);
endmodule

module UBCON_27_8 (O, I);
  output [27:8] O;
  input [27:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
  UB1DCON_11 U3 (O[11], I[11]);
  UB1DCON_12 U4 (O[12], I[12]);
  UB1DCON_13 U5 (O[13], I[13]);
  UB1DCON_14 U6 (O[14], I[14]);
  UB1DCON_15 U7 (O[15], I[15]);
  UB1DCON_16 U8 (O[16], I[16]);
  UB1DCON_17 U9 (O[17], I[17]);
  UB1DCON_18 U10 (O[18], I[18]);
  UB1DCON_19 U11 (O[19], I[19]);
  UB1DCON_20 U12 (O[20], I[20]);
  UB1DCON_21 U13 (O[21], I[21]);
  UB1DCON_22 U14 (O[22], I[22]);
  UB1DCON_23 U15 (O[23], I[23]);
  UB1DCON_24 U16 (O[24], I[24]);
  UB1DCON_25 U17 (O[25], I[25]);
  UB1DCON_26 U18 (O[26], I[26]);
  UB1DCON_27 U19 (O[27], I[27]);
endmodule

module UBCON_31_30 (O, I);
  output [31:30] O;
  input [31:30] I;
  UB1DCON_30 U0 (O[30], I[30]);
  UB1DCON_31 U1 (O[31], I[31]);
endmodule

module UBCON_33_32 (O, I);
  output [33:32] O;
  input [33:32] I;
  UB1DCON_32 U0 (O[32], I[32]);
  UB1DCON_33 U1 (O[33], I[33]);
endmodule

module UBCON_35_34 (O, I);
  output [35:34] O;
  input [35:34] I;
  UB1DCON_34 U0 (O[34], I[34]);
  UB1DCON_35 U1 (O[35], I[35]);
endmodule

module UBCON_39_38 (O, I);
  output [39:38] O;
  input [39:38] I;
  UB1DCON_38 U0 (O[38], I[38]);
  UB1DCON_39 U1 (O[39], I[39]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_3_2 (O, I);
  output [3:2] O;
  input [3:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
endmodule

module UBCON_41_40 (O, I);
  output [41:40] O;
  input [41:40] I;
  UB1DCON_40 U0 (O[40], I[40]);
  UB1DCON_41 U1 (O[41], I[41]);
endmodule

module UBCON_43_42 (O, I);
  output [43:42] O;
  input [43:42] I;
  UB1DCON_42 U0 (O[42], I[42]);
  UB1DCON_43 U1 (O[43], I[43]);
endmodule

module UBCON_47_46 (O, I);
  output [47:46] O;
  input [47:46] I;
  UB1DCON_46 U0 (O[46], I[46]);
  UB1DCON_47 U1 (O[47], I[47]);
endmodule

module UBCON_49_48 (O, I);
  output [49:48] O;
  input [49:48] I;
  UB1DCON_48 U0 (O[48], I[48]);
  UB1DCON_49 U1 (O[49], I[49]);
endmodule

module UBCON_51_50 (O, I);
  output [51:50] O;
  input [51:50] I;
  UB1DCON_50 U0 (O[50], I[50]);
  UB1DCON_51 U1 (O[51], I[51]);
endmodule

module UBCON_55_54 (O, I);
  output [55:54] O;
  input [55:54] I;
  UB1DCON_54 U0 (O[54], I[54]);
  UB1DCON_55 U1 (O[55], I[55]);
endmodule

module UBCON_57_56 (O, I);
  output [57:56] O;
  input [57:56] I;
  UB1DCON_56 U0 (O[56], I[56]);
  UB1DCON_57 U1 (O[57], I[57]);
endmodule

module UBCON_59_58 (O, I);
  output [59:58] O;
  input [59:58] I;
  UB1DCON_58 U0 (O[58], I[58]);
  UB1DCON_59 U1 (O[59], I[59]);
endmodule

module UBCON_63_62 (O, I);
  output [63:62] O;
  input [63:62] I;
  UB1DCON_62 U0 (O[62], I[62]);
  UB1DCON_63 U1 (O[63], I[63]);
endmodule

module UBCON_64_0 (O, I);
  output [64:0] O;
  input [64:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
  UB1DCON_28 U28 (O[28], I[28]);
  UB1DCON_29 U29 (O[29], I[29]);
  UB1DCON_30 U30 (O[30], I[30]);
  UB1DCON_31 U31 (O[31], I[31]);
  UB1DCON_32 U32 (O[32], I[32]);
  UB1DCON_33 U33 (O[33], I[33]);
  UB1DCON_34 U34 (O[34], I[34]);
  UB1DCON_35 U35 (O[35], I[35]);
  UB1DCON_36 U36 (O[36], I[36]);
  UB1DCON_37 U37 (O[37], I[37]);
  UB1DCON_38 U38 (O[38], I[38]);
  UB1DCON_39 U39 (O[39], I[39]);
  UB1DCON_40 U40 (O[40], I[40]);
  UB1DCON_41 U41 (O[41], I[41]);
  UB1DCON_42 U42 (O[42], I[42]);
  UB1DCON_43 U43 (O[43], I[43]);
  UB1DCON_44 U44 (O[44], I[44]);
  UB1DCON_45 U45 (O[45], I[45]);
  UB1DCON_46 U46 (O[46], I[46]);
  UB1DCON_47 U47 (O[47], I[47]);
  UB1DCON_48 U48 (O[48], I[48]);
  UB1DCON_49 U49 (O[49], I[49]);
  UB1DCON_50 U50 (O[50], I[50]);
  UB1DCON_51 U51 (O[51], I[51]);
  UB1DCON_52 U52 (O[52], I[52]);
  UB1DCON_53 U53 (O[53], I[53]);
  UB1DCON_54 U54 (O[54], I[54]);
  UB1DCON_55 U55 (O[55], I[55]);
  UB1DCON_56 U56 (O[56], I[56]);
  UB1DCON_57 U57 (O[57], I[57]);
  UB1DCON_58 U58 (O[58], I[58]);
  UB1DCON_59 U59 (O[59], I[59]);
  UB1DCON_60 U60 (O[60], I[60]);
  UB1DCON_61 U61 (O[61], I[61]);
  UB1DCON_62 U62 (O[62], I[62]);
  UB1DCON_63 U63 (O[63], I[63]);
  UB1DCON_64 U64 (O[64], I[64]);
endmodule

module UBCON_66_2 (O, I);
  output [66:2] O;
  input [66:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
  UB1DCON_9 U7 (O[9], I[9]);
  UB1DCON_10 U8 (O[10], I[10]);
  UB1DCON_11 U9 (O[11], I[11]);
  UB1DCON_12 U10 (O[12], I[12]);
  UB1DCON_13 U11 (O[13], I[13]);
  UB1DCON_14 U12 (O[14], I[14]);
  UB1DCON_15 U13 (O[15], I[15]);
  UB1DCON_16 U14 (O[16], I[16]);
  UB1DCON_17 U15 (O[17], I[17]);
  UB1DCON_18 U16 (O[18], I[18]);
  UB1DCON_19 U17 (O[19], I[19]);
  UB1DCON_20 U18 (O[20], I[20]);
  UB1DCON_21 U19 (O[21], I[21]);
  UB1DCON_22 U20 (O[22], I[22]);
  UB1DCON_23 U21 (O[23], I[23]);
  UB1DCON_24 U22 (O[24], I[24]);
  UB1DCON_25 U23 (O[25], I[25]);
  UB1DCON_26 U24 (O[26], I[26]);
  UB1DCON_27 U25 (O[27], I[27]);
  UB1DCON_28 U26 (O[28], I[28]);
  UB1DCON_29 U27 (O[29], I[29]);
  UB1DCON_30 U28 (O[30], I[30]);
  UB1DCON_31 U29 (O[31], I[31]);
  UB1DCON_32 U30 (O[32], I[32]);
  UB1DCON_33 U31 (O[33], I[33]);
  UB1DCON_34 U32 (O[34], I[34]);
  UB1DCON_35 U33 (O[35], I[35]);
  UB1DCON_36 U34 (O[36], I[36]);
  UB1DCON_37 U35 (O[37], I[37]);
  UB1DCON_38 U36 (O[38], I[38]);
  UB1DCON_39 U37 (O[39], I[39]);
  UB1DCON_40 U38 (O[40], I[40]);
  UB1DCON_41 U39 (O[41], I[41]);
  UB1DCON_42 U40 (O[42], I[42]);
  UB1DCON_43 U41 (O[43], I[43]);
  UB1DCON_44 U42 (O[44], I[44]);
  UB1DCON_45 U43 (O[45], I[45]);
  UB1DCON_46 U44 (O[46], I[46]);
  UB1DCON_47 U45 (O[47], I[47]);
  UB1DCON_48 U46 (O[48], I[48]);
  UB1DCON_49 U47 (O[49], I[49]);
  UB1DCON_50 U48 (O[50], I[50]);
  UB1DCON_51 U49 (O[51], I[51]);
  UB1DCON_52 U50 (O[52], I[52]);
  UB1DCON_53 U51 (O[53], I[53]);
  UB1DCON_54 U52 (O[54], I[54]);
  UB1DCON_55 U53 (O[55], I[55]);
  UB1DCON_56 U54 (O[56], I[56]);
  UB1DCON_57 U55 (O[57], I[57]);
  UB1DCON_58 U56 (O[58], I[58]);
  UB1DCON_59 U57 (O[59], I[59]);
  UB1DCON_60 U58 (O[60], I[60]);
  UB1DCON_61 U59 (O[61], I[61]);
  UB1DCON_62 U60 (O[62], I[62]);
  UB1DCON_63 U61 (O[63], I[63]);
  UB1DCON_64 U62 (O[64], I[64]);
  UB1DCON_65 U63 (O[65], I[65]);
  UB1DCON_66 U64 (O[66], I[66]);
endmodule

module UBCON_68_4 (O, I);
  output [68:4] O;
  input [68:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
  UB1DCON_19 U15 (O[19], I[19]);
  UB1DCON_20 U16 (O[20], I[20]);
  UB1DCON_21 U17 (O[21], I[21]);
  UB1DCON_22 U18 (O[22], I[22]);
  UB1DCON_23 U19 (O[23], I[23]);
  UB1DCON_24 U20 (O[24], I[24]);
  UB1DCON_25 U21 (O[25], I[25]);
  UB1DCON_26 U22 (O[26], I[26]);
  UB1DCON_27 U23 (O[27], I[27]);
  UB1DCON_28 U24 (O[28], I[28]);
  UB1DCON_29 U25 (O[29], I[29]);
  UB1DCON_30 U26 (O[30], I[30]);
  UB1DCON_31 U27 (O[31], I[31]);
  UB1DCON_32 U28 (O[32], I[32]);
  UB1DCON_33 U29 (O[33], I[33]);
  UB1DCON_34 U30 (O[34], I[34]);
  UB1DCON_35 U31 (O[35], I[35]);
  UB1DCON_36 U32 (O[36], I[36]);
  UB1DCON_37 U33 (O[37], I[37]);
  UB1DCON_38 U34 (O[38], I[38]);
  UB1DCON_39 U35 (O[39], I[39]);
  UB1DCON_40 U36 (O[40], I[40]);
  UB1DCON_41 U37 (O[41], I[41]);
  UB1DCON_42 U38 (O[42], I[42]);
  UB1DCON_43 U39 (O[43], I[43]);
  UB1DCON_44 U40 (O[44], I[44]);
  UB1DCON_45 U41 (O[45], I[45]);
  UB1DCON_46 U42 (O[46], I[46]);
  UB1DCON_47 U43 (O[47], I[47]);
  UB1DCON_48 U44 (O[48], I[48]);
  UB1DCON_49 U45 (O[49], I[49]);
  UB1DCON_50 U46 (O[50], I[50]);
  UB1DCON_51 U47 (O[51], I[51]);
  UB1DCON_52 U48 (O[52], I[52]);
  UB1DCON_53 U49 (O[53], I[53]);
  UB1DCON_54 U50 (O[54], I[54]);
  UB1DCON_55 U51 (O[55], I[55]);
  UB1DCON_56 U52 (O[56], I[56]);
  UB1DCON_57 U53 (O[57], I[57]);
  UB1DCON_58 U54 (O[58], I[58]);
  UB1DCON_59 U55 (O[59], I[59]);
  UB1DCON_60 U56 (O[60], I[60]);
  UB1DCON_61 U57 (O[61], I[61]);
  UB1DCON_62 U58 (O[62], I[62]);
  UB1DCON_63 U59 (O[63], I[63]);
  UB1DCON_64 U60 (O[64], I[64]);
  UB1DCON_65 U61 (O[65], I[65]);
  UB1DCON_66 U62 (O[66], I[66]);
  UB1DCON_67 U63 (O[67], I[67]);
  UB1DCON_68 U64 (O[68], I[68]);
endmodule

module UBCON_70_6 (O, I);
  output [70:6] O;
  input [70:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
  UB1DCON_9 U3 (O[9], I[9]);
  UB1DCON_10 U4 (O[10], I[10]);
  UB1DCON_11 U5 (O[11], I[11]);
  UB1DCON_12 U6 (O[12], I[12]);
  UB1DCON_13 U7 (O[13], I[13]);
  UB1DCON_14 U8 (O[14], I[14]);
  UB1DCON_15 U9 (O[15], I[15]);
  UB1DCON_16 U10 (O[16], I[16]);
  UB1DCON_17 U11 (O[17], I[17]);
  UB1DCON_18 U12 (O[18], I[18]);
  UB1DCON_19 U13 (O[19], I[19]);
  UB1DCON_20 U14 (O[20], I[20]);
  UB1DCON_21 U15 (O[21], I[21]);
  UB1DCON_22 U16 (O[22], I[22]);
  UB1DCON_23 U17 (O[23], I[23]);
  UB1DCON_24 U18 (O[24], I[24]);
  UB1DCON_25 U19 (O[25], I[25]);
  UB1DCON_26 U20 (O[26], I[26]);
  UB1DCON_27 U21 (O[27], I[27]);
  UB1DCON_28 U22 (O[28], I[28]);
  UB1DCON_29 U23 (O[29], I[29]);
  UB1DCON_30 U24 (O[30], I[30]);
  UB1DCON_31 U25 (O[31], I[31]);
  UB1DCON_32 U26 (O[32], I[32]);
  UB1DCON_33 U27 (O[33], I[33]);
  UB1DCON_34 U28 (O[34], I[34]);
  UB1DCON_35 U29 (O[35], I[35]);
  UB1DCON_36 U30 (O[36], I[36]);
  UB1DCON_37 U31 (O[37], I[37]);
  UB1DCON_38 U32 (O[38], I[38]);
  UB1DCON_39 U33 (O[39], I[39]);
  UB1DCON_40 U34 (O[40], I[40]);
  UB1DCON_41 U35 (O[41], I[41]);
  UB1DCON_42 U36 (O[42], I[42]);
  UB1DCON_43 U37 (O[43], I[43]);
  UB1DCON_44 U38 (O[44], I[44]);
  UB1DCON_45 U39 (O[45], I[45]);
  UB1DCON_46 U40 (O[46], I[46]);
  UB1DCON_47 U41 (O[47], I[47]);
  UB1DCON_48 U42 (O[48], I[48]);
  UB1DCON_49 U43 (O[49], I[49]);
  UB1DCON_50 U44 (O[50], I[50]);
  UB1DCON_51 U45 (O[51], I[51]);
  UB1DCON_52 U46 (O[52], I[52]);
  UB1DCON_53 U47 (O[53], I[53]);
  UB1DCON_54 U48 (O[54], I[54]);
  UB1DCON_55 U49 (O[55], I[55]);
  UB1DCON_56 U50 (O[56], I[56]);
  UB1DCON_57 U51 (O[57], I[57]);
  UB1DCON_58 U52 (O[58], I[58]);
  UB1DCON_59 U53 (O[59], I[59]);
  UB1DCON_60 U54 (O[60], I[60]);
  UB1DCON_61 U55 (O[61], I[61]);
  UB1DCON_62 U56 (O[62], I[62]);
  UB1DCON_63 U57 (O[63], I[63]);
  UB1DCON_64 U58 (O[64], I[64]);
  UB1DCON_65 U59 (O[65], I[65]);
  UB1DCON_66 U60 (O[66], I[66]);
  UB1DCON_67 U61 (O[67], I[67]);
  UB1DCON_68 U62 (O[68], I[68]);
  UB1DCON_69 U63 (O[69], I[69]);
  UB1DCON_70 U64 (O[70], I[70]);
endmodule

module UBCON_72_8 (O, I);
  output [72:8] O;
  input [72:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
  UB1DCON_11 U3 (O[11], I[11]);
  UB1DCON_12 U4 (O[12], I[12]);
  UB1DCON_13 U5 (O[13], I[13]);
  UB1DCON_14 U6 (O[14], I[14]);
  UB1DCON_15 U7 (O[15], I[15]);
  UB1DCON_16 U8 (O[16], I[16]);
  UB1DCON_17 U9 (O[17], I[17]);
  UB1DCON_18 U10 (O[18], I[18]);
  UB1DCON_19 U11 (O[19], I[19]);
  UB1DCON_20 U12 (O[20], I[20]);
  UB1DCON_21 U13 (O[21], I[21]);
  UB1DCON_22 U14 (O[22], I[22]);
  UB1DCON_23 U15 (O[23], I[23]);
  UB1DCON_24 U16 (O[24], I[24]);
  UB1DCON_25 U17 (O[25], I[25]);
  UB1DCON_26 U18 (O[26], I[26]);
  UB1DCON_27 U19 (O[27], I[27]);
  UB1DCON_28 U20 (O[28], I[28]);
  UB1DCON_29 U21 (O[29], I[29]);
  UB1DCON_30 U22 (O[30], I[30]);
  UB1DCON_31 U23 (O[31], I[31]);
  UB1DCON_32 U24 (O[32], I[32]);
  UB1DCON_33 U25 (O[33], I[33]);
  UB1DCON_34 U26 (O[34], I[34]);
  UB1DCON_35 U27 (O[35], I[35]);
  UB1DCON_36 U28 (O[36], I[36]);
  UB1DCON_37 U29 (O[37], I[37]);
  UB1DCON_38 U30 (O[38], I[38]);
  UB1DCON_39 U31 (O[39], I[39]);
  UB1DCON_40 U32 (O[40], I[40]);
  UB1DCON_41 U33 (O[41], I[41]);
  UB1DCON_42 U34 (O[42], I[42]);
  UB1DCON_43 U35 (O[43], I[43]);
  UB1DCON_44 U36 (O[44], I[44]);
  UB1DCON_45 U37 (O[45], I[45]);
  UB1DCON_46 U38 (O[46], I[46]);
  UB1DCON_47 U39 (O[47], I[47]);
  UB1DCON_48 U40 (O[48], I[48]);
  UB1DCON_49 U41 (O[49], I[49]);
  UB1DCON_50 U42 (O[50], I[50]);
  UB1DCON_51 U43 (O[51], I[51]);
  UB1DCON_52 U44 (O[52], I[52]);
  UB1DCON_53 U45 (O[53], I[53]);
  UB1DCON_54 U46 (O[54], I[54]);
  UB1DCON_55 U47 (O[55], I[55]);
  UB1DCON_56 U48 (O[56], I[56]);
  UB1DCON_57 U49 (O[57], I[57]);
  UB1DCON_58 U50 (O[58], I[58]);
  UB1DCON_59 U51 (O[59], I[59]);
  UB1DCON_60 U52 (O[60], I[60]);
  UB1DCON_61 U53 (O[61], I[61]);
  UB1DCON_62 U54 (O[62], I[62]);
  UB1DCON_63 U55 (O[63], I[63]);
  UB1DCON_64 U56 (O[64], I[64]);
  UB1DCON_65 U57 (O[65], I[65]);
  UB1DCON_66 U58 (O[66], I[66]);
  UB1DCON_67 U59 (O[67], I[67]);
  UB1DCON_68 U60 (O[68], I[68]);
  UB1DCON_69 U61 (O[69], I[69]);
  UB1DCON_70 U62 (O[70], I[70]);
  UB1DCON_71 U63 (O[71], I[71]);
  UB1DCON_72 U64 (O[72], I[72]);
endmodule

module UBCON_74_10 (O, I);
  output [74:10] O;
  input [74:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
  UB1DCON_13 U3 (O[13], I[13]);
  UB1DCON_14 U4 (O[14], I[14]);
  UB1DCON_15 U5 (O[15], I[15]);
  UB1DCON_16 U6 (O[16], I[16]);
  UB1DCON_17 U7 (O[17], I[17]);
  UB1DCON_18 U8 (O[18], I[18]);
  UB1DCON_19 U9 (O[19], I[19]);
  UB1DCON_20 U10 (O[20], I[20]);
  UB1DCON_21 U11 (O[21], I[21]);
  UB1DCON_22 U12 (O[22], I[22]);
  UB1DCON_23 U13 (O[23], I[23]);
  UB1DCON_24 U14 (O[24], I[24]);
  UB1DCON_25 U15 (O[25], I[25]);
  UB1DCON_26 U16 (O[26], I[26]);
  UB1DCON_27 U17 (O[27], I[27]);
  UB1DCON_28 U18 (O[28], I[28]);
  UB1DCON_29 U19 (O[29], I[29]);
  UB1DCON_30 U20 (O[30], I[30]);
  UB1DCON_31 U21 (O[31], I[31]);
  UB1DCON_32 U22 (O[32], I[32]);
  UB1DCON_33 U23 (O[33], I[33]);
  UB1DCON_34 U24 (O[34], I[34]);
  UB1DCON_35 U25 (O[35], I[35]);
  UB1DCON_36 U26 (O[36], I[36]);
  UB1DCON_37 U27 (O[37], I[37]);
  UB1DCON_38 U28 (O[38], I[38]);
  UB1DCON_39 U29 (O[39], I[39]);
  UB1DCON_40 U30 (O[40], I[40]);
  UB1DCON_41 U31 (O[41], I[41]);
  UB1DCON_42 U32 (O[42], I[42]);
  UB1DCON_43 U33 (O[43], I[43]);
  UB1DCON_44 U34 (O[44], I[44]);
  UB1DCON_45 U35 (O[45], I[45]);
  UB1DCON_46 U36 (O[46], I[46]);
  UB1DCON_47 U37 (O[47], I[47]);
  UB1DCON_48 U38 (O[48], I[48]);
  UB1DCON_49 U39 (O[49], I[49]);
  UB1DCON_50 U40 (O[50], I[50]);
  UB1DCON_51 U41 (O[51], I[51]);
  UB1DCON_52 U42 (O[52], I[52]);
  UB1DCON_53 U43 (O[53], I[53]);
  UB1DCON_54 U44 (O[54], I[54]);
  UB1DCON_55 U45 (O[55], I[55]);
  UB1DCON_56 U46 (O[56], I[56]);
  UB1DCON_57 U47 (O[57], I[57]);
  UB1DCON_58 U48 (O[58], I[58]);
  UB1DCON_59 U49 (O[59], I[59]);
  UB1DCON_60 U50 (O[60], I[60]);
  UB1DCON_61 U51 (O[61], I[61]);
  UB1DCON_62 U52 (O[62], I[62]);
  UB1DCON_63 U53 (O[63], I[63]);
  UB1DCON_64 U54 (O[64], I[64]);
  UB1DCON_65 U55 (O[65], I[65]);
  UB1DCON_66 U56 (O[66], I[66]);
  UB1DCON_67 U57 (O[67], I[67]);
  UB1DCON_68 U58 (O[68], I[68]);
  UB1DCON_69 U59 (O[69], I[69]);
  UB1DCON_70 U60 (O[70], I[70]);
  UB1DCON_71 U61 (O[71], I[71]);
  UB1DCON_72 U62 (O[72], I[72]);
  UB1DCON_73 U63 (O[73], I[73]);
  UB1DCON_74 U64 (O[74], I[74]);
endmodule

module UBCON_75_69 (O, I);
  output [75:69] O;
  input [75:69] I;
  UB1DCON_69 U0 (O[69], I[69]);
  UB1DCON_70 U1 (O[70], I[70]);
  UB1DCON_71 U2 (O[71], I[71]);
  UB1DCON_72 U3 (O[72], I[72]);
  UB1DCON_73 U4 (O[73], I[73]);
  UB1DCON_74 U5 (O[74], I[74]);
  UB1DCON_75 U6 (O[75], I[75]);
endmodule

module UBCON_76_12 (O, I);
  output [76:12] O;
  input [76:12] I;
  UB1DCON_12 U0 (O[12], I[12]);
  UB1DCON_13 U1 (O[13], I[13]);
  UB1DCON_14 U2 (O[14], I[14]);
  UB1DCON_15 U3 (O[15], I[15]);
  UB1DCON_16 U4 (O[16], I[16]);
  UB1DCON_17 U5 (O[17], I[17]);
  UB1DCON_18 U6 (O[18], I[18]);
  UB1DCON_19 U7 (O[19], I[19]);
  UB1DCON_20 U8 (O[20], I[20]);
  UB1DCON_21 U9 (O[21], I[21]);
  UB1DCON_22 U10 (O[22], I[22]);
  UB1DCON_23 U11 (O[23], I[23]);
  UB1DCON_24 U12 (O[24], I[24]);
  UB1DCON_25 U13 (O[25], I[25]);
  UB1DCON_26 U14 (O[26], I[26]);
  UB1DCON_27 U15 (O[27], I[27]);
  UB1DCON_28 U16 (O[28], I[28]);
  UB1DCON_29 U17 (O[29], I[29]);
  UB1DCON_30 U18 (O[30], I[30]);
  UB1DCON_31 U19 (O[31], I[31]);
  UB1DCON_32 U20 (O[32], I[32]);
  UB1DCON_33 U21 (O[33], I[33]);
  UB1DCON_34 U22 (O[34], I[34]);
  UB1DCON_35 U23 (O[35], I[35]);
  UB1DCON_36 U24 (O[36], I[36]);
  UB1DCON_37 U25 (O[37], I[37]);
  UB1DCON_38 U26 (O[38], I[38]);
  UB1DCON_39 U27 (O[39], I[39]);
  UB1DCON_40 U28 (O[40], I[40]);
  UB1DCON_41 U29 (O[41], I[41]);
  UB1DCON_42 U30 (O[42], I[42]);
  UB1DCON_43 U31 (O[43], I[43]);
  UB1DCON_44 U32 (O[44], I[44]);
  UB1DCON_45 U33 (O[45], I[45]);
  UB1DCON_46 U34 (O[46], I[46]);
  UB1DCON_47 U35 (O[47], I[47]);
  UB1DCON_48 U36 (O[48], I[48]);
  UB1DCON_49 U37 (O[49], I[49]);
  UB1DCON_50 U38 (O[50], I[50]);
  UB1DCON_51 U39 (O[51], I[51]);
  UB1DCON_52 U40 (O[52], I[52]);
  UB1DCON_53 U41 (O[53], I[53]);
  UB1DCON_54 U42 (O[54], I[54]);
  UB1DCON_55 U43 (O[55], I[55]);
  UB1DCON_56 U44 (O[56], I[56]);
  UB1DCON_57 U45 (O[57], I[57]);
  UB1DCON_58 U46 (O[58], I[58]);
  UB1DCON_59 U47 (O[59], I[59]);
  UB1DCON_60 U48 (O[60], I[60]);
  UB1DCON_61 U49 (O[61], I[61]);
  UB1DCON_62 U50 (O[62], I[62]);
  UB1DCON_63 U51 (O[63], I[63]);
  UB1DCON_64 U52 (O[64], I[64]);
  UB1DCON_65 U53 (O[65], I[65]);
  UB1DCON_66 U54 (O[66], I[66]);
  UB1DCON_67 U55 (O[67], I[67]);
  UB1DCON_68 U56 (O[68], I[68]);
  UB1DCON_69 U57 (O[69], I[69]);
  UB1DCON_70 U58 (O[70], I[70]);
  UB1DCON_71 U59 (O[71], I[71]);
  UB1DCON_72 U60 (O[72], I[72]);
  UB1DCON_73 U61 (O[73], I[73]);
  UB1DCON_74 U62 (O[74], I[74]);
  UB1DCON_75 U63 (O[75], I[75]);
  UB1DCON_76 U64 (O[76], I[76]);
endmodule

module UBCON_78_14 (O, I);
  output [78:14] O;
  input [78:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
  UB1DCON_18 U4 (O[18], I[18]);
  UB1DCON_19 U5 (O[19], I[19]);
  UB1DCON_20 U6 (O[20], I[20]);
  UB1DCON_21 U7 (O[21], I[21]);
  UB1DCON_22 U8 (O[22], I[22]);
  UB1DCON_23 U9 (O[23], I[23]);
  UB1DCON_24 U10 (O[24], I[24]);
  UB1DCON_25 U11 (O[25], I[25]);
  UB1DCON_26 U12 (O[26], I[26]);
  UB1DCON_27 U13 (O[27], I[27]);
  UB1DCON_28 U14 (O[28], I[28]);
  UB1DCON_29 U15 (O[29], I[29]);
  UB1DCON_30 U16 (O[30], I[30]);
  UB1DCON_31 U17 (O[31], I[31]);
  UB1DCON_32 U18 (O[32], I[32]);
  UB1DCON_33 U19 (O[33], I[33]);
  UB1DCON_34 U20 (O[34], I[34]);
  UB1DCON_35 U21 (O[35], I[35]);
  UB1DCON_36 U22 (O[36], I[36]);
  UB1DCON_37 U23 (O[37], I[37]);
  UB1DCON_38 U24 (O[38], I[38]);
  UB1DCON_39 U25 (O[39], I[39]);
  UB1DCON_40 U26 (O[40], I[40]);
  UB1DCON_41 U27 (O[41], I[41]);
  UB1DCON_42 U28 (O[42], I[42]);
  UB1DCON_43 U29 (O[43], I[43]);
  UB1DCON_44 U30 (O[44], I[44]);
  UB1DCON_45 U31 (O[45], I[45]);
  UB1DCON_46 U32 (O[46], I[46]);
  UB1DCON_47 U33 (O[47], I[47]);
  UB1DCON_48 U34 (O[48], I[48]);
  UB1DCON_49 U35 (O[49], I[49]);
  UB1DCON_50 U36 (O[50], I[50]);
  UB1DCON_51 U37 (O[51], I[51]);
  UB1DCON_52 U38 (O[52], I[52]);
  UB1DCON_53 U39 (O[53], I[53]);
  UB1DCON_54 U40 (O[54], I[54]);
  UB1DCON_55 U41 (O[55], I[55]);
  UB1DCON_56 U42 (O[56], I[56]);
  UB1DCON_57 U43 (O[57], I[57]);
  UB1DCON_58 U44 (O[58], I[58]);
  UB1DCON_59 U45 (O[59], I[59]);
  UB1DCON_60 U46 (O[60], I[60]);
  UB1DCON_61 U47 (O[61], I[61]);
  UB1DCON_62 U48 (O[62], I[62]);
  UB1DCON_63 U49 (O[63], I[63]);
  UB1DCON_64 U50 (O[64], I[64]);
  UB1DCON_65 U51 (O[65], I[65]);
  UB1DCON_66 U52 (O[66], I[66]);
  UB1DCON_67 U53 (O[67], I[67]);
  UB1DCON_68 U54 (O[68], I[68]);
  UB1DCON_69 U55 (O[69], I[69]);
  UB1DCON_70 U56 (O[70], I[70]);
  UB1DCON_71 U57 (O[71], I[71]);
  UB1DCON_72 U58 (O[72], I[72]);
  UB1DCON_73 U59 (O[73], I[73]);
  UB1DCON_74 U60 (O[74], I[74]);
  UB1DCON_75 U61 (O[75], I[75]);
  UB1DCON_76 U62 (O[76], I[76]);
  UB1DCON_77 U63 (O[77], I[77]);
  UB1DCON_78 U64 (O[78], I[78]);
endmodule

module UBCON_7_6 (O, I);
  output [7:6] O;
  input [7:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
endmodule

module UBCON_80_16 (O, I);
  output [80:16] O;
  input [80:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
  UB1DCON_19 U3 (O[19], I[19]);
  UB1DCON_20 U4 (O[20], I[20]);
  UB1DCON_21 U5 (O[21], I[21]);
  UB1DCON_22 U6 (O[22], I[22]);
  UB1DCON_23 U7 (O[23], I[23]);
  UB1DCON_24 U8 (O[24], I[24]);
  UB1DCON_25 U9 (O[25], I[25]);
  UB1DCON_26 U10 (O[26], I[26]);
  UB1DCON_27 U11 (O[27], I[27]);
  UB1DCON_28 U12 (O[28], I[28]);
  UB1DCON_29 U13 (O[29], I[29]);
  UB1DCON_30 U14 (O[30], I[30]);
  UB1DCON_31 U15 (O[31], I[31]);
  UB1DCON_32 U16 (O[32], I[32]);
  UB1DCON_33 U17 (O[33], I[33]);
  UB1DCON_34 U18 (O[34], I[34]);
  UB1DCON_35 U19 (O[35], I[35]);
  UB1DCON_36 U20 (O[36], I[36]);
  UB1DCON_37 U21 (O[37], I[37]);
  UB1DCON_38 U22 (O[38], I[38]);
  UB1DCON_39 U23 (O[39], I[39]);
  UB1DCON_40 U24 (O[40], I[40]);
  UB1DCON_41 U25 (O[41], I[41]);
  UB1DCON_42 U26 (O[42], I[42]);
  UB1DCON_43 U27 (O[43], I[43]);
  UB1DCON_44 U28 (O[44], I[44]);
  UB1DCON_45 U29 (O[45], I[45]);
  UB1DCON_46 U30 (O[46], I[46]);
  UB1DCON_47 U31 (O[47], I[47]);
  UB1DCON_48 U32 (O[48], I[48]);
  UB1DCON_49 U33 (O[49], I[49]);
  UB1DCON_50 U34 (O[50], I[50]);
  UB1DCON_51 U35 (O[51], I[51]);
  UB1DCON_52 U36 (O[52], I[52]);
  UB1DCON_53 U37 (O[53], I[53]);
  UB1DCON_54 U38 (O[54], I[54]);
  UB1DCON_55 U39 (O[55], I[55]);
  UB1DCON_56 U40 (O[56], I[56]);
  UB1DCON_57 U41 (O[57], I[57]);
  UB1DCON_58 U42 (O[58], I[58]);
  UB1DCON_59 U43 (O[59], I[59]);
  UB1DCON_60 U44 (O[60], I[60]);
  UB1DCON_61 U45 (O[61], I[61]);
  UB1DCON_62 U46 (O[62], I[62]);
  UB1DCON_63 U47 (O[63], I[63]);
  UB1DCON_64 U48 (O[64], I[64]);
  UB1DCON_65 U49 (O[65], I[65]);
  UB1DCON_66 U50 (O[66], I[66]);
  UB1DCON_67 U51 (O[67], I[67]);
  UB1DCON_68 U52 (O[68], I[68]);
  UB1DCON_69 U53 (O[69], I[69]);
  UB1DCON_70 U54 (O[70], I[70]);
  UB1DCON_71 U55 (O[71], I[71]);
  UB1DCON_72 U56 (O[72], I[72]);
  UB1DCON_73 U57 (O[73], I[73]);
  UB1DCON_74 U58 (O[74], I[74]);
  UB1DCON_75 U59 (O[75], I[75]);
  UB1DCON_76 U60 (O[76], I[76]);
  UB1DCON_77 U61 (O[77], I[77]);
  UB1DCON_78 U62 (O[78], I[78]);
  UB1DCON_79 U63 (O[79], I[79]);
  UB1DCON_80 U64 (O[80], I[80]);
endmodule

module UBCON_82_18 (O, I);
  output [82:18] O;
  input [82:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
  UB1DCON_20 U2 (O[20], I[20]);
  UB1DCON_21 U3 (O[21], I[21]);
  UB1DCON_22 U4 (O[22], I[22]);
  UB1DCON_23 U5 (O[23], I[23]);
  UB1DCON_24 U6 (O[24], I[24]);
  UB1DCON_25 U7 (O[25], I[25]);
  UB1DCON_26 U8 (O[26], I[26]);
  UB1DCON_27 U9 (O[27], I[27]);
  UB1DCON_28 U10 (O[28], I[28]);
  UB1DCON_29 U11 (O[29], I[29]);
  UB1DCON_30 U12 (O[30], I[30]);
  UB1DCON_31 U13 (O[31], I[31]);
  UB1DCON_32 U14 (O[32], I[32]);
  UB1DCON_33 U15 (O[33], I[33]);
  UB1DCON_34 U16 (O[34], I[34]);
  UB1DCON_35 U17 (O[35], I[35]);
  UB1DCON_36 U18 (O[36], I[36]);
  UB1DCON_37 U19 (O[37], I[37]);
  UB1DCON_38 U20 (O[38], I[38]);
  UB1DCON_39 U21 (O[39], I[39]);
  UB1DCON_40 U22 (O[40], I[40]);
  UB1DCON_41 U23 (O[41], I[41]);
  UB1DCON_42 U24 (O[42], I[42]);
  UB1DCON_43 U25 (O[43], I[43]);
  UB1DCON_44 U26 (O[44], I[44]);
  UB1DCON_45 U27 (O[45], I[45]);
  UB1DCON_46 U28 (O[46], I[46]);
  UB1DCON_47 U29 (O[47], I[47]);
  UB1DCON_48 U30 (O[48], I[48]);
  UB1DCON_49 U31 (O[49], I[49]);
  UB1DCON_50 U32 (O[50], I[50]);
  UB1DCON_51 U33 (O[51], I[51]);
  UB1DCON_52 U34 (O[52], I[52]);
  UB1DCON_53 U35 (O[53], I[53]);
  UB1DCON_54 U36 (O[54], I[54]);
  UB1DCON_55 U37 (O[55], I[55]);
  UB1DCON_56 U38 (O[56], I[56]);
  UB1DCON_57 U39 (O[57], I[57]);
  UB1DCON_58 U40 (O[58], I[58]);
  UB1DCON_59 U41 (O[59], I[59]);
  UB1DCON_60 U42 (O[60], I[60]);
  UB1DCON_61 U43 (O[61], I[61]);
  UB1DCON_62 U44 (O[62], I[62]);
  UB1DCON_63 U45 (O[63], I[63]);
  UB1DCON_64 U46 (O[64], I[64]);
  UB1DCON_65 U47 (O[65], I[65]);
  UB1DCON_66 U48 (O[66], I[66]);
  UB1DCON_67 U49 (O[67], I[67]);
  UB1DCON_68 U50 (O[68], I[68]);
  UB1DCON_69 U51 (O[69], I[69]);
  UB1DCON_70 U52 (O[70], I[70]);
  UB1DCON_71 U53 (O[71], I[71]);
  UB1DCON_72 U54 (O[72], I[72]);
  UB1DCON_73 U55 (O[73], I[73]);
  UB1DCON_74 U56 (O[74], I[74]);
  UB1DCON_75 U57 (O[75], I[75]);
  UB1DCON_76 U58 (O[76], I[76]);
  UB1DCON_77 U59 (O[77], I[77]);
  UB1DCON_78 U60 (O[78], I[78]);
  UB1DCON_79 U61 (O[79], I[79]);
  UB1DCON_80 U62 (O[80], I[80]);
  UB1DCON_81 U63 (O[81], I[81]);
  UB1DCON_82 U64 (O[82], I[82]);
endmodule

module UBCON_83_77 (O, I);
  output [83:77] O;
  input [83:77] I;
  UB1DCON_77 U0 (O[77], I[77]);
  UB1DCON_78 U1 (O[78], I[78]);
  UB1DCON_79 U2 (O[79], I[79]);
  UB1DCON_80 U3 (O[80], I[80]);
  UB1DCON_81 U4 (O[81], I[81]);
  UB1DCON_82 U5 (O[82], I[82]);
  UB1DCON_83 U6 (O[83], I[83]);
endmodule

module UBCON_84_20 (O, I);
  output [84:20] O;
  input [84:20] I;
  UB1DCON_20 U0 (O[20], I[20]);
  UB1DCON_21 U1 (O[21], I[21]);
  UB1DCON_22 U2 (O[22], I[22]);
  UB1DCON_23 U3 (O[23], I[23]);
  UB1DCON_24 U4 (O[24], I[24]);
  UB1DCON_25 U5 (O[25], I[25]);
  UB1DCON_26 U6 (O[26], I[26]);
  UB1DCON_27 U7 (O[27], I[27]);
  UB1DCON_28 U8 (O[28], I[28]);
  UB1DCON_29 U9 (O[29], I[29]);
  UB1DCON_30 U10 (O[30], I[30]);
  UB1DCON_31 U11 (O[31], I[31]);
  UB1DCON_32 U12 (O[32], I[32]);
  UB1DCON_33 U13 (O[33], I[33]);
  UB1DCON_34 U14 (O[34], I[34]);
  UB1DCON_35 U15 (O[35], I[35]);
  UB1DCON_36 U16 (O[36], I[36]);
  UB1DCON_37 U17 (O[37], I[37]);
  UB1DCON_38 U18 (O[38], I[38]);
  UB1DCON_39 U19 (O[39], I[39]);
  UB1DCON_40 U20 (O[40], I[40]);
  UB1DCON_41 U21 (O[41], I[41]);
  UB1DCON_42 U22 (O[42], I[42]);
  UB1DCON_43 U23 (O[43], I[43]);
  UB1DCON_44 U24 (O[44], I[44]);
  UB1DCON_45 U25 (O[45], I[45]);
  UB1DCON_46 U26 (O[46], I[46]);
  UB1DCON_47 U27 (O[47], I[47]);
  UB1DCON_48 U28 (O[48], I[48]);
  UB1DCON_49 U29 (O[49], I[49]);
  UB1DCON_50 U30 (O[50], I[50]);
  UB1DCON_51 U31 (O[51], I[51]);
  UB1DCON_52 U32 (O[52], I[52]);
  UB1DCON_53 U33 (O[53], I[53]);
  UB1DCON_54 U34 (O[54], I[54]);
  UB1DCON_55 U35 (O[55], I[55]);
  UB1DCON_56 U36 (O[56], I[56]);
  UB1DCON_57 U37 (O[57], I[57]);
  UB1DCON_58 U38 (O[58], I[58]);
  UB1DCON_59 U39 (O[59], I[59]);
  UB1DCON_60 U40 (O[60], I[60]);
  UB1DCON_61 U41 (O[61], I[61]);
  UB1DCON_62 U42 (O[62], I[62]);
  UB1DCON_63 U43 (O[63], I[63]);
  UB1DCON_64 U44 (O[64], I[64]);
  UB1DCON_65 U45 (O[65], I[65]);
  UB1DCON_66 U46 (O[66], I[66]);
  UB1DCON_67 U47 (O[67], I[67]);
  UB1DCON_68 U48 (O[68], I[68]);
  UB1DCON_69 U49 (O[69], I[69]);
  UB1DCON_70 U50 (O[70], I[70]);
  UB1DCON_71 U51 (O[71], I[71]);
  UB1DCON_72 U52 (O[72], I[72]);
  UB1DCON_73 U53 (O[73], I[73]);
  UB1DCON_74 U54 (O[74], I[74]);
  UB1DCON_75 U55 (O[75], I[75]);
  UB1DCON_76 U56 (O[76], I[76]);
  UB1DCON_77 U57 (O[77], I[77]);
  UB1DCON_78 U58 (O[78], I[78]);
  UB1DCON_79 U59 (O[79], I[79]);
  UB1DCON_80 U60 (O[80], I[80]);
  UB1DCON_81 U61 (O[81], I[81]);
  UB1DCON_82 U62 (O[82], I[82]);
  UB1DCON_83 U63 (O[83], I[83]);
  UB1DCON_84 U64 (O[84], I[84]);
endmodule

module UBCON_86_22 (O, I);
  output [86:22] O;
  input [86:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
  UB1DCON_24 U2 (O[24], I[24]);
  UB1DCON_25 U3 (O[25], I[25]);
  UB1DCON_26 U4 (O[26], I[26]);
  UB1DCON_27 U5 (O[27], I[27]);
  UB1DCON_28 U6 (O[28], I[28]);
  UB1DCON_29 U7 (O[29], I[29]);
  UB1DCON_30 U8 (O[30], I[30]);
  UB1DCON_31 U9 (O[31], I[31]);
  UB1DCON_32 U10 (O[32], I[32]);
  UB1DCON_33 U11 (O[33], I[33]);
  UB1DCON_34 U12 (O[34], I[34]);
  UB1DCON_35 U13 (O[35], I[35]);
  UB1DCON_36 U14 (O[36], I[36]);
  UB1DCON_37 U15 (O[37], I[37]);
  UB1DCON_38 U16 (O[38], I[38]);
  UB1DCON_39 U17 (O[39], I[39]);
  UB1DCON_40 U18 (O[40], I[40]);
  UB1DCON_41 U19 (O[41], I[41]);
  UB1DCON_42 U20 (O[42], I[42]);
  UB1DCON_43 U21 (O[43], I[43]);
  UB1DCON_44 U22 (O[44], I[44]);
  UB1DCON_45 U23 (O[45], I[45]);
  UB1DCON_46 U24 (O[46], I[46]);
  UB1DCON_47 U25 (O[47], I[47]);
  UB1DCON_48 U26 (O[48], I[48]);
  UB1DCON_49 U27 (O[49], I[49]);
  UB1DCON_50 U28 (O[50], I[50]);
  UB1DCON_51 U29 (O[51], I[51]);
  UB1DCON_52 U30 (O[52], I[52]);
  UB1DCON_53 U31 (O[53], I[53]);
  UB1DCON_54 U32 (O[54], I[54]);
  UB1DCON_55 U33 (O[55], I[55]);
  UB1DCON_56 U34 (O[56], I[56]);
  UB1DCON_57 U35 (O[57], I[57]);
  UB1DCON_58 U36 (O[58], I[58]);
  UB1DCON_59 U37 (O[59], I[59]);
  UB1DCON_60 U38 (O[60], I[60]);
  UB1DCON_61 U39 (O[61], I[61]);
  UB1DCON_62 U40 (O[62], I[62]);
  UB1DCON_63 U41 (O[63], I[63]);
  UB1DCON_64 U42 (O[64], I[64]);
  UB1DCON_65 U43 (O[65], I[65]);
  UB1DCON_66 U44 (O[66], I[66]);
  UB1DCON_67 U45 (O[67], I[67]);
  UB1DCON_68 U46 (O[68], I[68]);
  UB1DCON_69 U47 (O[69], I[69]);
  UB1DCON_70 U48 (O[70], I[70]);
  UB1DCON_71 U49 (O[71], I[71]);
  UB1DCON_72 U50 (O[72], I[72]);
  UB1DCON_73 U51 (O[73], I[73]);
  UB1DCON_74 U52 (O[74], I[74]);
  UB1DCON_75 U53 (O[75], I[75]);
  UB1DCON_76 U54 (O[76], I[76]);
  UB1DCON_77 U55 (O[77], I[77]);
  UB1DCON_78 U56 (O[78], I[78]);
  UB1DCON_79 U57 (O[79], I[79]);
  UB1DCON_80 U58 (O[80], I[80]);
  UB1DCON_81 U59 (O[81], I[81]);
  UB1DCON_82 U60 (O[82], I[82]);
  UB1DCON_83 U61 (O[83], I[83]);
  UB1DCON_84 U62 (O[84], I[84]);
  UB1DCON_85 U63 (O[85], I[85]);
  UB1DCON_86 U64 (O[86], I[86]);
endmodule

module UBCON_88_24 (O, I);
  output [88:24] O;
  input [88:24] I;
  UB1DCON_24 U0 (O[24], I[24]);
  UB1DCON_25 U1 (O[25], I[25]);
  UB1DCON_26 U2 (O[26], I[26]);
  UB1DCON_27 U3 (O[27], I[27]);
  UB1DCON_28 U4 (O[28], I[28]);
  UB1DCON_29 U5 (O[29], I[29]);
  UB1DCON_30 U6 (O[30], I[30]);
  UB1DCON_31 U7 (O[31], I[31]);
  UB1DCON_32 U8 (O[32], I[32]);
  UB1DCON_33 U9 (O[33], I[33]);
  UB1DCON_34 U10 (O[34], I[34]);
  UB1DCON_35 U11 (O[35], I[35]);
  UB1DCON_36 U12 (O[36], I[36]);
  UB1DCON_37 U13 (O[37], I[37]);
  UB1DCON_38 U14 (O[38], I[38]);
  UB1DCON_39 U15 (O[39], I[39]);
  UB1DCON_40 U16 (O[40], I[40]);
  UB1DCON_41 U17 (O[41], I[41]);
  UB1DCON_42 U18 (O[42], I[42]);
  UB1DCON_43 U19 (O[43], I[43]);
  UB1DCON_44 U20 (O[44], I[44]);
  UB1DCON_45 U21 (O[45], I[45]);
  UB1DCON_46 U22 (O[46], I[46]);
  UB1DCON_47 U23 (O[47], I[47]);
  UB1DCON_48 U24 (O[48], I[48]);
  UB1DCON_49 U25 (O[49], I[49]);
  UB1DCON_50 U26 (O[50], I[50]);
  UB1DCON_51 U27 (O[51], I[51]);
  UB1DCON_52 U28 (O[52], I[52]);
  UB1DCON_53 U29 (O[53], I[53]);
  UB1DCON_54 U30 (O[54], I[54]);
  UB1DCON_55 U31 (O[55], I[55]);
  UB1DCON_56 U32 (O[56], I[56]);
  UB1DCON_57 U33 (O[57], I[57]);
  UB1DCON_58 U34 (O[58], I[58]);
  UB1DCON_59 U35 (O[59], I[59]);
  UB1DCON_60 U36 (O[60], I[60]);
  UB1DCON_61 U37 (O[61], I[61]);
  UB1DCON_62 U38 (O[62], I[62]);
  UB1DCON_63 U39 (O[63], I[63]);
  UB1DCON_64 U40 (O[64], I[64]);
  UB1DCON_65 U41 (O[65], I[65]);
  UB1DCON_66 U42 (O[66], I[66]);
  UB1DCON_67 U43 (O[67], I[67]);
  UB1DCON_68 U44 (O[68], I[68]);
  UB1DCON_69 U45 (O[69], I[69]);
  UB1DCON_70 U46 (O[70], I[70]);
  UB1DCON_71 U47 (O[71], I[71]);
  UB1DCON_72 U48 (O[72], I[72]);
  UB1DCON_73 U49 (O[73], I[73]);
  UB1DCON_74 U50 (O[74], I[74]);
  UB1DCON_75 U51 (O[75], I[75]);
  UB1DCON_76 U52 (O[76], I[76]);
  UB1DCON_77 U53 (O[77], I[77]);
  UB1DCON_78 U54 (O[78], I[78]);
  UB1DCON_79 U55 (O[79], I[79]);
  UB1DCON_80 U56 (O[80], I[80]);
  UB1DCON_81 U57 (O[81], I[81]);
  UB1DCON_82 U58 (O[82], I[82]);
  UB1DCON_83 U59 (O[83], I[83]);
  UB1DCON_84 U60 (O[84], I[84]);
  UB1DCON_85 U61 (O[85], I[85]);
  UB1DCON_86 U62 (O[86], I[86]);
  UB1DCON_87 U63 (O[87], I[87]);
  UB1DCON_88 U64 (O[88], I[88]);
endmodule

module UBCON_90_26 (O, I);
  output [90:26] O;
  input [90:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
  UB1DCON_28 U2 (O[28], I[28]);
  UB1DCON_29 U3 (O[29], I[29]);
  UB1DCON_30 U4 (O[30], I[30]);
  UB1DCON_31 U5 (O[31], I[31]);
  UB1DCON_32 U6 (O[32], I[32]);
  UB1DCON_33 U7 (O[33], I[33]);
  UB1DCON_34 U8 (O[34], I[34]);
  UB1DCON_35 U9 (O[35], I[35]);
  UB1DCON_36 U10 (O[36], I[36]);
  UB1DCON_37 U11 (O[37], I[37]);
  UB1DCON_38 U12 (O[38], I[38]);
  UB1DCON_39 U13 (O[39], I[39]);
  UB1DCON_40 U14 (O[40], I[40]);
  UB1DCON_41 U15 (O[41], I[41]);
  UB1DCON_42 U16 (O[42], I[42]);
  UB1DCON_43 U17 (O[43], I[43]);
  UB1DCON_44 U18 (O[44], I[44]);
  UB1DCON_45 U19 (O[45], I[45]);
  UB1DCON_46 U20 (O[46], I[46]);
  UB1DCON_47 U21 (O[47], I[47]);
  UB1DCON_48 U22 (O[48], I[48]);
  UB1DCON_49 U23 (O[49], I[49]);
  UB1DCON_50 U24 (O[50], I[50]);
  UB1DCON_51 U25 (O[51], I[51]);
  UB1DCON_52 U26 (O[52], I[52]);
  UB1DCON_53 U27 (O[53], I[53]);
  UB1DCON_54 U28 (O[54], I[54]);
  UB1DCON_55 U29 (O[55], I[55]);
  UB1DCON_56 U30 (O[56], I[56]);
  UB1DCON_57 U31 (O[57], I[57]);
  UB1DCON_58 U32 (O[58], I[58]);
  UB1DCON_59 U33 (O[59], I[59]);
  UB1DCON_60 U34 (O[60], I[60]);
  UB1DCON_61 U35 (O[61], I[61]);
  UB1DCON_62 U36 (O[62], I[62]);
  UB1DCON_63 U37 (O[63], I[63]);
  UB1DCON_64 U38 (O[64], I[64]);
  UB1DCON_65 U39 (O[65], I[65]);
  UB1DCON_66 U40 (O[66], I[66]);
  UB1DCON_67 U41 (O[67], I[67]);
  UB1DCON_68 U42 (O[68], I[68]);
  UB1DCON_69 U43 (O[69], I[69]);
  UB1DCON_70 U44 (O[70], I[70]);
  UB1DCON_71 U45 (O[71], I[71]);
  UB1DCON_72 U46 (O[72], I[72]);
  UB1DCON_73 U47 (O[73], I[73]);
  UB1DCON_74 U48 (O[74], I[74]);
  UB1DCON_75 U49 (O[75], I[75]);
  UB1DCON_76 U50 (O[76], I[76]);
  UB1DCON_77 U51 (O[77], I[77]);
  UB1DCON_78 U52 (O[78], I[78]);
  UB1DCON_79 U53 (O[79], I[79]);
  UB1DCON_80 U54 (O[80], I[80]);
  UB1DCON_81 U55 (O[81], I[81]);
  UB1DCON_82 U56 (O[82], I[82]);
  UB1DCON_83 U57 (O[83], I[83]);
  UB1DCON_84 U58 (O[84], I[84]);
  UB1DCON_85 U59 (O[85], I[85]);
  UB1DCON_86 U60 (O[86], I[86]);
  UB1DCON_87 U61 (O[87], I[87]);
  UB1DCON_88 U62 (O[88], I[88]);
  UB1DCON_89 U63 (O[89], I[89]);
  UB1DCON_90 U64 (O[90], I[90]);
endmodule

module UBCON_91_85 (O, I);
  output [91:85] O;
  input [91:85] I;
  UB1DCON_85 U0 (O[85], I[85]);
  UB1DCON_86 U1 (O[86], I[86]);
  UB1DCON_87 U2 (O[87], I[87]);
  UB1DCON_88 U3 (O[88], I[88]);
  UB1DCON_89 U4 (O[89], I[89]);
  UB1DCON_90 U5 (O[90], I[90]);
  UB1DCON_91 U6 (O[91], I[91]);
endmodule

module UBCON_92_28 (O, I);
  output [92:28] O;
  input [92:28] I;
  UB1DCON_28 U0 (O[28], I[28]);
  UB1DCON_29 U1 (O[29], I[29]);
  UB1DCON_30 U2 (O[30], I[30]);
  UB1DCON_31 U3 (O[31], I[31]);
  UB1DCON_32 U4 (O[32], I[32]);
  UB1DCON_33 U5 (O[33], I[33]);
  UB1DCON_34 U6 (O[34], I[34]);
  UB1DCON_35 U7 (O[35], I[35]);
  UB1DCON_36 U8 (O[36], I[36]);
  UB1DCON_37 U9 (O[37], I[37]);
  UB1DCON_38 U10 (O[38], I[38]);
  UB1DCON_39 U11 (O[39], I[39]);
  UB1DCON_40 U12 (O[40], I[40]);
  UB1DCON_41 U13 (O[41], I[41]);
  UB1DCON_42 U14 (O[42], I[42]);
  UB1DCON_43 U15 (O[43], I[43]);
  UB1DCON_44 U16 (O[44], I[44]);
  UB1DCON_45 U17 (O[45], I[45]);
  UB1DCON_46 U18 (O[46], I[46]);
  UB1DCON_47 U19 (O[47], I[47]);
  UB1DCON_48 U20 (O[48], I[48]);
  UB1DCON_49 U21 (O[49], I[49]);
  UB1DCON_50 U22 (O[50], I[50]);
  UB1DCON_51 U23 (O[51], I[51]);
  UB1DCON_52 U24 (O[52], I[52]);
  UB1DCON_53 U25 (O[53], I[53]);
  UB1DCON_54 U26 (O[54], I[54]);
  UB1DCON_55 U27 (O[55], I[55]);
  UB1DCON_56 U28 (O[56], I[56]);
  UB1DCON_57 U29 (O[57], I[57]);
  UB1DCON_58 U30 (O[58], I[58]);
  UB1DCON_59 U31 (O[59], I[59]);
  UB1DCON_60 U32 (O[60], I[60]);
  UB1DCON_61 U33 (O[61], I[61]);
  UB1DCON_62 U34 (O[62], I[62]);
  UB1DCON_63 U35 (O[63], I[63]);
  UB1DCON_64 U36 (O[64], I[64]);
  UB1DCON_65 U37 (O[65], I[65]);
  UB1DCON_66 U38 (O[66], I[66]);
  UB1DCON_67 U39 (O[67], I[67]);
  UB1DCON_68 U40 (O[68], I[68]);
  UB1DCON_69 U41 (O[69], I[69]);
  UB1DCON_70 U42 (O[70], I[70]);
  UB1DCON_71 U43 (O[71], I[71]);
  UB1DCON_72 U44 (O[72], I[72]);
  UB1DCON_73 U45 (O[73], I[73]);
  UB1DCON_74 U46 (O[74], I[74]);
  UB1DCON_75 U47 (O[75], I[75]);
  UB1DCON_76 U48 (O[76], I[76]);
  UB1DCON_77 U49 (O[77], I[77]);
  UB1DCON_78 U50 (O[78], I[78]);
  UB1DCON_79 U51 (O[79], I[79]);
  UB1DCON_80 U52 (O[80], I[80]);
  UB1DCON_81 U53 (O[81], I[81]);
  UB1DCON_82 U54 (O[82], I[82]);
  UB1DCON_83 U55 (O[83], I[83]);
  UB1DCON_84 U56 (O[84], I[84]);
  UB1DCON_85 U57 (O[85], I[85]);
  UB1DCON_86 U58 (O[86], I[86]);
  UB1DCON_87 U59 (O[87], I[87]);
  UB1DCON_88 U60 (O[88], I[88]);
  UB1DCON_89 U61 (O[89], I[89]);
  UB1DCON_90 U62 (O[90], I[90]);
  UB1DCON_91 U63 (O[91], I[91]);
  UB1DCON_92 U64 (O[92], I[92]);
endmodule

module UBCON_94_30 (O, I);
  output [94:30] O;
  input [94:30] I;
  UB1DCON_30 U0 (O[30], I[30]);
  UB1DCON_31 U1 (O[31], I[31]);
  UB1DCON_32 U2 (O[32], I[32]);
  UB1DCON_33 U3 (O[33], I[33]);
  UB1DCON_34 U4 (O[34], I[34]);
  UB1DCON_35 U5 (O[35], I[35]);
  UB1DCON_36 U6 (O[36], I[36]);
  UB1DCON_37 U7 (O[37], I[37]);
  UB1DCON_38 U8 (O[38], I[38]);
  UB1DCON_39 U9 (O[39], I[39]);
  UB1DCON_40 U10 (O[40], I[40]);
  UB1DCON_41 U11 (O[41], I[41]);
  UB1DCON_42 U12 (O[42], I[42]);
  UB1DCON_43 U13 (O[43], I[43]);
  UB1DCON_44 U14 (O[44], I[44]);
  UB1DCON_45 U15 (O[45], I[45]);
  UB1DCON_46 U16 (O[46], I[46]);
  UB1DCON_47 U17 (O[47], I[47]);
  UB1DCON_48 U18 (O[48], I[48]);
  UB1DCON_49 U19 (O[49], I[49]);
  UB1DCON_50 U20 (O[50], I[50]);
  UB1DCON_51 U21 (O[51], I[51]);
  UB1DCON_52 U22 (O[52], I[52]);
  UB1DCON_53 U23 (O[53], I[53]);
  UB1DCON_54 U24 (O[54], I[54]);
  UB1DCON_55 U25 (O[55], I[55]);
  UB1DCON_56 U26 (O[56], I[56]);
  UB1DCON_57 U27 (O[57], I[57]);
  UB1DCON_58 U28 (O[58], I[58]);
  UB1DCON_59 U29 (O[59], I[59]);
  UB1DCON_60 U30 (O[60], I[60]);
  UB1DCON_61 U31 (O[61], I[61]);
  UB1DCON_62 U32 (O[62], I[62]);
  UB1DCON_63 U33 (O[63], I[63]);
  UB1DCON_64 U34 (O[64], I[64]);
  UB1DCON_65 U35 (O[65], I[65]);
  UB1DCON_66 U36 (O[66], I[66]);
  UB1DCON_67 U37 (O[67], I[67]);
  UB1DCON_68 U38 (O[68], I[68]);
  UB1DCON_69 U39 (O[69], I[69]);
  UB1DCON_70 U40 (O[70], I[70]);
  UB1DCON_71 U41 (O[71], I[71]);
  UB1DCON_72 U42 (O[72], I[72]);
  UB1DCON_73 U43 (O[73], I[73]);
  UB1DCON_74 U44 (O[74], I[74]);
  UB1DCON_75 U45 (O[75], I[75]);
  UB1DCON_76 U46 (O[76], I[76]);
  UB1DCON_77 U47 (O[77], I[77]);
  UB1DCON_78 U48 (O[78], I[78]);
  UB1DCON_79 U49 (O[79], I[79]);
  UB1DCON_80 U50 (O[80], I[80]);
  UB1DCON_81 U51 (O[81], I[81]);
  UB1DCON_82 U52 (O[82], I[82]);
  UB1DCON_83 U53 (O[83], I[83]);
  UB1DCON_84 U54 (O[84], I[84]);
  UB1DCON_85 U55 (O[85], I[85]);
  UB1DCON_86 U56 (O[86], I[86]);
  UB1DCON_87 U57 (O[87], I[87]);
  UB1DCON_88 U58 (O[88], I[88]);
  UB1DCON_89 U59 (O[89], I[89]);
  UB1DCON_90 U60 (O[90], I[90]);
  UB1DCON_91 U61 (O[91], I[91]);
  UB1DCON_92 U62 (O[92], I[92]);
  UB1DCON_93 U63 (O[93], I[93]);
  UB1DCON_94 U64 (O[94], I[94]);
endmodule

module UBCON_96_32 (O, I);
  output [96:32] O;
  input [96:32] I;
  UB1DCON_32 U0 (O[32], I[32]);
  UB1DCON_33 U1 (O[33], I[33]);
  UB1DCON_34 U2 (O[34], I[34]);
  UB1DCON_35 U3 (O[35], I[35]);
  UB1DCON_36 U4 (O[36], I[36]);
  UB1DCON_37 U5 (O[37], I[37]);
  UB1DCON_38 U6 (O[38], I[38]);
  UB1DCON_39 U7 (O[39], I[39]);
  UB1DCON_40 U8 (O[40], I[40]);
  UB1DCON_41 U9 (O[41], I[41]);
  UB1DCON_42 U10 (O[42], I[42]);
  UB1DCON_43 U11 (O[43], I[43]);
  UB1DCON_44 U12 (O[44], I[44]);
  UB1DCON_45 U13 (O[45], I[45]);
  UB1DCON_46 U14 (O[46], I[46]);
  UB1DCON_47 U15 (O[47], I[47]);
  UB1DCON_48 U16 (O[48], I[48]);
  UB1DCON_49 U17 (O[49], I[49]);
  UB1DCON_50 U18 (O[50], I[50]);
  UB1DCON_51 U19 (O[51], I[51]);
  UB1DCON_52 U20 (O[52], I[52]);
  UB1DCON_53 U21 (O[53], I[53]);
  UB1DCON_54 U22 (O[54], I[54]);
  UB1DCON_55 U23 (O[55], I[55]);
  UB1DCON_56 U24 (O[56], I[56]);
  UB1DCON_57 U25 (O[57], I[57]);
  UB1DCON_58 U26 (O[58], I[58]);
  UB1DCON_59 U27 (O[59], I[59]);
  UB1DCON_60 U28 (O[60], I[60]);
  UB1DCON_61 U29 (O[61], I[61]);
  UB1DCON_62 U30 (O[62], I[62]);
  UB1DCON_63 U31 (O[63], I[63]);
  UB1DCON_64 U32 (O[64], I[64]);
  UB1DCON_65 U33 (O[65], I[65]);
  UB1DCON_66 U34 (O[66], I[66]);
  UB1DCON_67 U35 (O[67], I[67]);
  UB1DCON_68 U36 (O[68], I[68]);
  UB1DCON_69 U37 (O[69], I[69]);
  UB1DCON_70 U38 (O[70], I[70]);
  UB1DCON_71 U39 (O[71], I[71]);
  UB1DCON_72 U40 (O[72], I[72]);
  UB1DCON_73 U41 (O[73], I[73]);
  UB1DCON_74 U42 (O[74], I[74]);
  UB1DCON_75 U43 (O[75], I[75]);
  UB1DCON_76 U44 (O[76], I[76]);
  UB1DCON_77 U45 (O[77], I[77]);
  UB1DCON_78 U46 (O[78], I[78]);
  UB1DCON_79 U47 (O[79], I[79]);
  UB1DCON_80 U48 (O[80], I[80]);
  UB1DCON_81 U49 (O[81], I[81]);
  UB1DCON_82 U50 (O[82], I[82]);
  UB1DCON_83 U51 (O[83], I[83]);
  UB1DCON_84 U52 (O[84], I[84]);
  UB1DCON_85 U53 (O[85], I[85]);
  UB1DCON_86 U54 (O[86], I[86]);
  UB1DCON_87 U55 (O[87], I[87]);
  UB1DCON_88 U56 (O[88], I[88]);
  UB1DCON_89 U57 (O[89], I[89]);
  UB1DCON_90 U58 (O[90], I[90]);
  UB1DCON_91 U59 (O[91], I[91]);
  UB1DCON_92 U60 (O[92], I[92]);
  UB1DCON_93 U61 (O[93], I[93]);
  UB1DCON_94 U62 (O[94], I[94]);
  UB1DCON_95 U63 (O[95], I[95]);
  UB1DCON_96 U64 (O[96], I[96]);
endmodule

module UBCON_98_34 (O, I);
  output [98:34] O;
  input [98:34] I;
  UB1DCON_34 U0 (O[34], I[34]);
  UB1DCON_35 U1 (O[35], I[35]);
  UB1DCON_36 U2 (O[36], I[36]);
  UB1DCON_37 U3 (O[37], I[37]);
  UB1DCON_38 U4 (O[38], I[38]);
  UB1DCON_39 U5 (O[39], I[39]);
  UB1DCON_40 U6 (O[40], I[40]);
  UB1DCON_41 U7 (O[41], I[41]);
  UB1DCON_42 U8 (O[42], I[42]);
  UB1DCON_43 U9 (O[43], I[43]);
  UB1DCON_44 U10 (O[44], I[44]);
  UB1DCON_45 U11 (O[45], I[45]);
  UB1DCON_46 U12 (O[46], I[46]);
  UB1DCON_47 U13 (O[47], I[47]);
  UB1DCON_48 U14 (O[48], I[48]);
  UB1DCON_49 U15 (O[49], I[49]);
  UB1DCON_50 U16 (O[50], I[50]);
  UB1DCON_51 U17 (O[51], I[51]);
  UB1DCON_52 U18 (O[52], I[52]);
  UB1DCON_53 U19 (O[53], I[53]);
  UB1DCON_54 U20 (O[54], I[54]);
  UB1DCON_55 U21 (O[55], I[55]);
  UB1DCON_56 U22 (O[56], I[56]);
  UB1DCON_57 U23 (O[57], I[57]);
  UB1DCON_58 U24 (O[58], I[58]);
  UB1DCON_59 U25 (O[59], I[59]);
  UB1DCON_60 U26 (O[60], I[60]);
  UB1DCON_61 U27 (O[61], I[61]);
  UB1DCON_62 U28 (O[62], I[62]);
  UB1DCON_63 U29 (O[63], I[63]);
  UB1DCON_64 U30 (O[64], I[64]);
  UB1DCON_65 U31 (O[65], I[65]);
  UB1DCON_66 U32 (O[66], I[66]);
  UB1DCON_67 U33 (O[67], I[67]);
  UB1DCON_68 U34 (O[68], I[68]);
  UB1DCON_69 U35 (O[69], I[69]);
  UB1DCON_70 U36 (O[70], I[70]);
  UB1DCON_71 U37 (O[71], I[71]);
  UB1DCON_72 U38 (O[72], I[72]);
  UB1DCON_73 U39 (O[73], I[73]);
  UB1DCON_74 U40 (O[74], I[74]);
  UB1DCON_75 U41 (O[75], I[75]);
  UB1DCON_76 U42 (O[76], I[76]);
  UB1DCON_77 U43 (O[77], I[77]);
  UB1DCON_78 U44 (O[78], I[78]);
  UB1DCON_79 U45 (O[79], I[79]);
  UB1DCON_80 U46 (O[80], I[80]);
  UB1DCON_81 U47 (O[81], I[81]);
  UB1DCON_82 U48 (O[82], I[82]);
  UB1DCON_83 U49 (O[83], I[83]);
  UB1DCON_84 U50 (O[84], I[84]);
  UB1DCON_85 U51 (O[85], I[85]);
  UB1DCON_86 U52 (O[86], I[86]);
  UB1DCON_87 U53 (O[87], I[87]);
  UB1DCON_88 U54 (O[88], I[88]);
  UB1DCON_89 U55 (O[89], I[89]);
  UB1DCON_90 U56 (O[90], I[90]);
  UB1DCON_91 U57 (O[91], I[91]);
  UB1DCON_92 U58 (O[92], I[92]);
  UB1DCON_93 U59 (O[93], I[93]);
  UB1DCON_94 U60 (O[94], I[94]);
  UB1DCON_95 U61 (O[95], I[95]);
  UB1DCON_96 U62 (O[96], I[96]);
  UB1DCON_97 U63 (O[97], I[97]);
  UB1DCON_98 U64 (O[98], I[98]);
endmodule

module UBCON_99_93 (O, I);
  output [99:93] O;
  input [99:93] I;
  UB1DCON_93 U0 (O[93], I[93]);
  UB1DCON_94 U1 (O[94], I[94]);
  UB1DCON_95 U2 (O[95], I[95]);
  UB1DCON_96 U3 (O[96], I[96]);
  UB1DCON_97 U4 (O[97], I[97]);
  UB1DCON_98 U5 (O[98], I[98]);
  UB1DCON_99 U6 (O[99], I[99]);
endmodule

module UBCSe_126_0_126_0 (S, X, Y);
  output [127:0] S;
  input [126:0] X;
  input [126:0] Y;
  UBPureCSe_126_0 U0 (S[127:0], X[126:0], Y[126:0]);
endmodule

module UBPureCSe_126_0 (S, X, Y);
  output [127:0] S;
  input [126:0] X;
  input [126:0] Y;
  wire C;
  UBPriCSlA_126_0 U0 (S, X, Y, C);
  UBZero_0_0 U1 (C);
endmodule

module UBRCB_0_0 (Co, S, X, Y, Ci);
  output Co;
  output S;
  input Ci;
  input X;
  input Y;
  UBFA_0 U0 (Co, S, X, Y, Ci);
endmodule

module UBRCB_105_92 (Co, S, X, Y, Ci);
  output Co;
  output [105:92] S;
  input Ci;
  input [105:92] X;
  input [105:92] Y;
  wire C100;
  wire C101;
  wire C102;
  wire C103;
  wire C104;
  wire C105;
  wire C93;
  wire C94;
  wire C95;
  wire C96;
  wire C97;
  wire C98;
  wire C99;
  UBFA_92 U0 (C93, S[92], X[92], Y[92], Ci);
  UBFA_93 U1 (C94, S[93], X[93], Y[93], C93);
  UBFA_94 U2 (C95, S[94], X[94], Y[94], C94);
  UBFA_95 U3 (C96, S[95], X[95], Y[95], C95);
  UBFA_96 U4 (C97, S[96], X[96], Y[96], C96);
  UBFA_97 U5 (C98, S[97], X[97], Y[97], C97);
  UBFA_98 U6 (C99, S[98], X[98], Y[98], C98);
  UBFA_99 U7 (C100, S[99], X[99], Y[99], C99);
  UBFA_100 U8 (C101, S[100], X[100], Y[100], C100);
  UBFA_101 U9 (C102, S[101], X[101], Y[101], C101);
  UBFA_102 U10 (C103, S[102], X[102], Y[102], C102);
  UBFA_103 U11 (C104, S[103], X[103], Y[103], C103);
  UBFA_104 U12 (C105, S[104], X[104], Y[104], C104);
  UBFA_105 U13 (Co, S[105], X[105], Y[105], C105);
endmodule

module UBRCB_10_7 (Co, S, X, Y, Ci);
  output Co;
  output [10:7] S;
  input Ci;
  input [10:7] X;
  input [10:7] Y;
  wire C10;
  wire C8;
  wire C9;
  UBFA_7 U0 (C8, S[7], X[7], Y[7], Ci);
  UBFA_8 U1 (C9, S[8], X[8], Y[8], C8);
  UBFA_9 U2 (C10, S[9], X[9], Y[9], C9);
  UBFA_10 U3 (Co, S[10], X[10], Y[10], C10);
endmodule

module UBRCB_120_106 (Co, S, X, Y, Ci);
  output Co;
  output [120:106] S;
  input Ci;
  input [120:106] X;
  input [120:106] Y;
  wire C107;
  wire C108;
  wire C109;
  wire C110;
  wire C111;
  wire C112;
  wire C113;
  wire C114;
  wire C115;
  wire C116;
  wire C117;
  wire C118;
  wire C119;
  wire C120;
  UBFA_106 U0 (C107, S[106], X[106], Y[106], Ci);
  UBFA_107 U1 (C108, S[107], X[107], Y[107], C107);
  UBFA_108 U2 (C109, S[108], X[108], Y[108], C108);
  UBFA_109 U3 (C110, S[109], X[109], Y[109], C109);
  UBFA_110 U4 (C111, S[110], X[110], Y[110], C110);
  UBFA_111 U5 (C112, S[111], X[111], Y[111], C111);
  UBFA_112 U6 (C113, S[112], X[112], Y[112], C112);
  UBFA_113 U7 (C114, S[113], X[113], Y[113], C113);
  UBFA_114 U8 (C115, S[114], X[114], Y[114], C114);
  UBFA_115 U9 (C116, S[115], X[115], Y[115], C115);
  UBFA_116 U10 (C117, S[116], X[116], Y[116], C116);
  UBFA_117 U11 (C118, S[117], X[117], Y[117], C117);
  UBFA_118 U12 (C119, S[118], X[118], Y[118], C118);
  UBFA_119 U13 (C120, S[119], X[119], Y[119], C119);
  UBFA_120 U14 (Co, S[120], X[120], Y[120], C120);
endmodule

module UBRCB_126_121 (Co, S, X, Y, Ci);
  output Co;
  output [126:121] S;
  input Ci;
  input [126:121] X;
  input [126:121] Y;
  wire C122;
  wire C123;
  wire C124;
  wire C125;
  wire C126;
  UBFA_121 U0 (C122, S[121], X[121], Y[121], Ci);
  UBFA_122 U1 (C123, S[122], X[122], Y[122], C122);
  UBFA_123 U2 (C124, S[123], X[123], Y[123], C123);
  UBFA_124 U3 (C125, S[124], X[124], Y[124], C124);
  UBFA_125 U4 (C126, S[125], X[125], Y[125], C125);
  UBFA_126 U5 (Co, S[126], X[126], Y[126], C126);
endmodule

module UBRCB_15_11 (Co, S, X, Y, Ci);
  output Co;
  output [15:11] S;
  input Ci;
  input [15:11] X;
  input [15:11] Y;
  wire C12;
  wire C13;
  wire C14;
  wire C15;
  UBFA_11 U0 (C12, S[11], X[11], Y[11], Ci);
  UBFA_12 U1 (C13, S[12], X[12], Y[12], C12);
  UBFA_13 U2 (C14, S[13], X[13], Y[13], C13);
  UBFA_14 U3 (C15, S[14], X[14], Y[14], C14);
  UBFA_15 U4 (Co, S[15], X[15], Y[15], C15);
endmodule

module UBRCB_1_1 (Co, S, X, Y, Ci);
  output Co;
  output S;
  input Ci;
  input X;
  input Y;
  UBFA_1 U0 (Co, S, X, Y, Ci);
endmodule

module UBRCB_21_16 (Co, S, X, Y, Ci);
  output Co;
  output [21:16] S;
  input Ci;
  input [21:16] X;
  input [21:16] Y;
  wire C17;
  wire C18;
  wire C19;
  wire C20;
  wire C21;
  UBFA_16 U0 (C17, S[16], X[16], Y[16], Ci);
  UBFA_17 U1 (C18, S[17], X[17], Y[17], C17);
  UBFA_18 U2 (C19, S[18], X[18], Y[18], C18);
  UBFA_19 U3 (C20, S[19], X[19], Y[19], C19);
  UBFA_20 U4 (C21, S[20], X[20], Y[20], C20);
  UBFA_21 U5 (Co, S[21], X[21], Y[21], C21);
endmodule

module UBRCB_28_22 (Co, S, X, Y, Ci);
  output Co;
  output [28:22] S;
  input Ci;
  input [28:22] X;
  input [28:22] Y;
  wire C23;
  wire C24;
  wire C25;
  wire C26;
  wire C27;
  wire C28;
  UBFA_22 U0 (C23, S[22], X[22], Y[22], Ci);
  UBFA_23 U1 (C24, S[23], X[23], Y[23], C23);
  UBFA_24 U2 (C25, S[24], X[24], Y[24], C24);
  UBFA_25 U3 (C26, S[25], X[25], Y[25], C25);
  UBFA_26 U4 (C27, S[26], X[26], Y[26], C26);
  UBFA_27 U5 (C28, S[27], X[27], Y[27], C27);
  UBFA_28 U6 (Co, S[28], X[28], Y[28], C28);
endmodule

module UBRCB_36_29 (Co, S, X, Y, Ci);
  output Co;
  output [36:29] S;
  input Ci;
  input [36:29] X;
  input [36:29] Y;
  wire C30;
  wire C31;
  wire C32;
  wire C33;
  wire C34;
  wire C35;
  wire C36;
  UBFA_29 U0 (C30, S[29], X[29], Y[29], Ci);
  UBFA_30 U1 (C31, S[30], X[30], Y[30], C30);
  UBFA_31 U2 (C32, S[31], X[31], Y[31], C31);
  UBFA_32 U3 (C33, S[32], X[32], Y[32], C32);
  UBFA_33 U4 (C34, S[33], X[33], Y[33], C33);
  UBFA_34 U5 (C35, S[34], X[34], Y[34], C34);
  UBFA_35 U6 (C36, S[35], X[35], Y[35], C35);
  UBFA_36 U7 (Co, S[36], X[36], Y[36], C36);
endmodule

module UBRCB_3_2 (Co, S, X, Y, Ci);
  output Co;
  output [3:2] S;
  input Ci;
  input [3:2] X;
  input [3:2] Y;
  wire C3;
  UBFA_2 U0 (C3, S[2], X[2], Y[2], Ci);
  UBFA_3 U1 (Co, S[3], X[3], Y[3], C3);
endmodule

module UBRCB_45_37 (Co, S, X, Y, Ci);
  output Co;
  output [45:37] S;
  input Ci;
  input [45:37] X;
  input [45:37] Y;
  wire C38;
  wire C39;
  wire C40;
  wire C41;
  wire C42;
  wire C43;
  wire C44;
  wire C45;
  UBFA_37 U0 (C38, S[37], X[37], Y[37], Ci);
  UBFA_38 U1 (C39, S[38], X[38], Y[38], C38);
  UBFA_39 U2 (C40, S[39], X[39], Y[39], C39);
  UBFA_40 U3 (C41, S[40], X[40], Y[40], C40);
  UBFA_41 U4 (C42, S[41], X[41], Y[41], C41);
  UBFA_42 U5 (C43, S[42], X[42], Y[42], C42);
  UBFA_43 U6 (C44, S[43], X[43], Y[43], C43);
  UBFA_44 U7 (C45, S[44], X[44], Y[44], C44);
  UBFA_45 U8 (Co, S[45], X[45], Y[45], C45);
endmodule

module UBRCB_55_46 (Co, S, X, Y, Ci);
  output Co;
  output [55:46] S;
  input Ci;
  input [55:46] X;
  input [55:46] Y;
  wire C47;
  wire C48;
  wire C49;
  wire C50;
  wire C51;
  wire C52;
  wire C53;
  wire C54;
  wire C55;
  UBFA_46 U0 (C47, S[46], X[46], Y[46], Ci);
  UBFA_47 U1 (C48, S[47], X[47], Y[47], C47);
  UBFA_48 U2 (C49, S[48], X[48], Y[48], C48);
  UBFA_49 U3 (C50, S[49], X[49], Y[49], C49);
  UBFA_50 U4 (C51, S[50], X[50], Y[50], C50);
  UBFA_51 U5 (C52, S[51], X[51], Y[51], C51);
  UBFA_52 U6 (C53, S[52], X[52], Y[52], C52);
  UBFA_53 U7 (C54, S[53], X[53], Y[53], C53);
  UBFA_54 U8 (C55, S[54], X[54], Y[54], C54);
  UBFA_55 U9 (Co, S[55], X[55], Y[55], C55);
endmodule

module UBRCB_66_56 (Co, S, X, Y, Ci);
  output Co;
  output [66:56] S;
  input Ci;
  input [66:56] X;
  input [66:56] Y;
  wire C57;
  wire C58;
  wire C59;
  wire C60;
  wire C61;
  wire C62;
  wire C63;
  wire C64;
  wire C65;
  wire C66;
  UBFA_56 U0 (C57, S[56], X[56], Y[56], Ci);
  UBFA_57 U1 (C58, S[57], X[57], Y[57], C57);
  UBFA_58 U2 (C59, S[58], X[58], Y[58], C58);
  UBFA_59 U3 (C60, S[59], X[59], Y[59], C59);
  UBFA_60 U4 (C61, S[60], X[60], Y[60], C60);
  UBFA_61 U5 (C62, S[61], X[61], Y[61], C61);
  UBFA_62 U6 (C63, S[62], X[62], Y[62], C62);
  UBFA_63 U7 (C64, S[63], X[63], Y[63], C63);
  UBFA_64 U8 (C65, S[64], X[64], Y[64], C64);
  UBFA_65 U9 (C66, S[65], X[65], Y[65], C65);
  UBFA_66 U10 (Co, S[66], X[66], Y[66], C66);
endmodule

module UBRCB_6_4 (Co, S, X, Y, Ci);
  output Co;
  output [6:4] S;
  input Ci;
  input [6:4] X;
  input [6:4] Y;
  wire C5;
  wire C6;
  UBFA_4 U0 (C5, S[4], X[4], Y[4], Ci);
  UBFA_5 U1 (C6, S[5], X[5], Y[5], C5);
  UBFA_6 U2 (Co, S[6], X[6], Y[6], C6);
endmodule

module UBRCB_78_67 (Co, S, X, Y, Ci);
  output Co;
  output [78:67] S;
  input Ci;
  input [78:67] X;
  input [78:67] Y;
  wire C68;
  wire C69;
  wire C70;
  wire C71;
  wire C72;
  wire C73;
  wire C74;
  wire C75;
  wire C76;
  wire C77;
  wire C78;
  UBFA_67 U0 (C68, S[67], X[67], Y[67], Ci);
  UBFA_68 U1 (C69, S[68], X[68], Y[68], C68);
  UBFA_69 U2 (C70, S[69], X[69], Y[69], C69);
  UBFA_70 U3 (C71, S[70], X[70], Y[70], C70);
  UBFA_71 U4 (C72, S[71], X[71], Y[71], C71);
  UBFA_72 U5 (C73, S[72], X[72], Y[72], C72);
  UBFA_73 U6 (C74, S[73], X[73], Y[73], C73);
  UBFA_74 U7 (C75, S[74], X[74], Y[74], C74);
  UBFA_75 U8 (C76, S[75], X[75], Y[75], C75);
  UBFA_76 U9 (C77, S[76], X[76], Y[76], C76);
  UBFA_77 U10 (C78, S[77], X[77], Y[77], C77);
  UBFA_78 U11 (Co, S[78], X[78], Y[78], C78);
endmodule

module UBRCB_91_79 (Co, S, X, Y, Ci);
  output Co;
  output [91:79] S;
  input Ci;
  input [91:79] X;
  input [91:79] Y;
  wire C80;
  wire C81;
  wire C82;
  wire C83;
  wire C84;
  wire C85;
  wire C86;
  wire C87;
  wire C88;
  wire C89;
  wire C90;
  wire C91;
  UBFA_79 U0 (C80, S[79], X[79], Y[79], Ci);
  UBFA_80 U1 (C81, S[80], X[80], Y[80], C80);
  UBFA_81 U2 (C82, S[81], X[81], Y[81], C81);
  UBFA_82 U3 (C83, S[82], X[82], Y[82], C82);
  UBFA_83 U4 (C84, S[83], X[83], Y[83], C83);
  UBFA_84 U5 (C85, S[84], X[84], Y[84], C84);
  UBFA_85 U6 (C86, S[85], X[85], Y[85], C85);
  UBFA_86 U7 (C87, S[86], X[86], Y[86], C86);
  UBFA_87 U8 (C88, S[87], X[87], Y[87], C87);
  UBFA_88 U9 (C89, S[88], X[88], Y[88], C88);
  UBFA_89 U10 (C90, S[89], X[89], Y[89], C89);
  UBFA_90 U11 (C91, S[90], X[90], Y[90], C90);
  UBFA_91 U12 (Co, S[91], X[91], Y[91], C91);
endmodule

module UBTCCONV127_127_0 (O, I);
  output [127:0] O;
  input [127:0] I;
  UBTC1CON127_0 U0 (O[0], I[0]);
  UBTC1CON127_1 U1 (O[1], I[1]);
  UBTC1CON127_2 U2 (O[2], I[2]);
  UBTC1CON127_3 U3 (O[3], I[3]);
  UBTC1CON127_4 U4 (O[4], I[4]);
  UBTC1CON127_5 U5 (O[5], I[5]);
  UBTC1CON127_6 U6 (O[6], I[6]);
  UBTC1CON127_7 U7 (O[7], I[7]);
  UBTC1CON127_8 U8 (O[8], I[8]);
  UBTC1CON127_9 U9 (O[9], I[9]);
  UBTC1CON127_10 U10 (O[10], I[10]);
  UBTC1CON127_11 U11 (O[11], I[11]);
  UBTC1CON127_12 U12 (O[12], I[12]);
  UBTC1CON127_13 U13 (O[13], I[13]);
  UBTC1CON127_14 U14 (O[14], I[14]);
  UBTC1CON127_15 U15 (O[15], I[15]);
  UBTC1CON127_16 U16 (O[16], I[16]);
  UBTC1CON127_17 U17 (O[17], I[17]);
  UBTC1CON127_18 U18 (O[18], I[18]);
  UBTC1CON127_19 U19 (O[19], I[19]);
  UBTC1CON127_20 U20 (O[20], I[20]);
  UBTC1CON127_21 U21 (O[21], I[21]);
  UBTC1CON127_22 U22 (O[22], I[22]);
  UBTC1CON127_23 U23 (O[23], I[23]);
  UBTC1CON127_24 U24 (O[24], I[24]);
  UBTC1CON127_25 U25 (O[25], I[25]);
  UBTC1CON127_26 U26 (O[26], I[26]);
  UBTC1CON127_27 U27 (O[27], I[27]);
  UBTC1CON127_28 U28 (O[28], I[28]);
  UBTC1CON127_29 U29 (O[29], I[29]);
  UBTC1CON127_30 U30 (O[30], I[30]);
  UBTC1CON127_31 U31 (O[31], I[31]);
  UBTC1CON127_32 U32 (O[32], I[32]);
  UBTC1CON127_33 U33 (O[33], I[33]);
  UBTC1CON127_34 U34 (O[34], I[34]);
  UBTC1CON127_35 U35 (O[35], I[35]);
  UBTC1CON127_36 U36 (O[36], I[36]);
  UBTC1CON127_37 U37 (O[37], I[37]);
  UBTC1CON127_38 U38 (O[38], I[38]);
  UBTC1CON127_39 U39 (O[39], I[39]);
  UBTC1CON127_40 U40 (O[40], I[40]);
  UBTC1CON127_41 U41 (O[41], I[41]);
  UBTC1CON127_42 U42 (O[42], I[42]);
  UBTC1CON127_43 U43 (O[43], I[43]);
  UBTC1CON127_44 U44 (O[44], I[44]);
  UBTC1CON127_45 U45 (O[45], I[45]);
  UBTC1CON127_46 U46 (O[46], I[46]);
  UBTC1CON127_47 U47 (O[47], I[47]);
  UBTC1CON127_48 U48 (O[48], I[48]);
  UBTC1CON127_49 U49 (O[49], I[49]);
  UBTC1CON127_50 U50 (O[50], I[50]);
  UBTC1CON127_51 U51 (O[51], I[51]);
  UBTC1CON127_52 U52 (O[52], I[52]);
  UBTC1CON127_53 U53 (O[53], I[53]);
  UBTC1CON127_54 U54 (O[54], I[54]);
  UBTC1CON127_55 U55 (O[55], I[55]);
  UBTC1CON127_56 U56 (O[56], I[56]);
  UBTC1CON127_57 U57 (O[57], I[57]);
  UBTC1CON127_58 U58 (O[58], I[58]);
  UBTC1CON127_59 U59 (O[59], I[59]);
  UBTC1CON127_60 U60 (O[60], I[60]);
  UBTC1CON127_61 U61 (O[61], I[61]);
  UBTC1CON127_62 U62 (O[62], I[62]);
  UBTC1CON127_63 U63 (O[63], I[63]);
  UBTC1CON127_64 U64 (O[64], I[64]);
  UBTC1CON127_65 U65 (O[65], I[65]);
  UBTC1CON127_66 U66 (O[66], I[66]);
  UBTC1CON127_67 U67 (O[67], I[67]);
  UBTC1CON127_68 U68 (O[68], I[68]);
  UBTC1CON127_69 U69 (O[69], I[69]);
  UBTC1CON127_70 U70 (O[70], I[70]);
  UBTC1CON127_71 U71 (O[71], I[71]);
  UBTC1CON127_72 U72 (O[72], I[72]);
  UBTC1CON127_73 U73 (O[73], I[73]);
  UBTC1CON127_74 U74 (O[74], I[74]);
  UBTC1CON127_75 U75 (O[75], I[75]);
  UBTC1CON127_76 U76 (O[76], I[76]);
  UBTC1CON127_77 U77 (O[77], I[77]);
  UBTC1CON127_78 U78 (O[78], I[78]);
  UBTC1CON127_79 U79 (O[79], I[79]);
  UBTC1CON127_80 U80 (O[80], I[80]);
  UBTC1CON127_81 U81 (O[81], I[81]);
  UBTC1CON127_82 U82 (O[82], I[82]);
  UBTC1CON127_83 U83 (O[83], I[83]);
  UBTC1CON127_84 U84 (O[84], I[84]);
  UBTC1CON127_85 U85 (O[85], I[85]);
  UBTC1CON127_86 U86 (O[86], I[86]);
  UBTC1CON127_87 U87 (O[87], I[87]);
  UBTC1CON127_88 U88 (O[88], I[88]);
  UBTC1CON127_89 U89 (O[89], I[89]);
  UBTC1CON127_90 U90 (O[90], I[90]);
  UBTC1CON127_91 U91 (O[91], I[91]);
  UBTC1CON127_92 U92 (O[92], I[92]);
  UBTC1CON127_93 U93 (O[93], I[93]);
  UBTC1CON127_94 U94 (O[94], I[94]);
  UBTC1CON127_95 U95 (O[95], I[95]);
  UBTC1CON127_96 U96 (O[96], I[96]);
  UBTC1CON127_97 U97 (O[97], I[97]);
  UBTC1CON127_98 U98 (O[98], I[98]);
  UBTC1CON127_99 U99 (O[99], I[99]);
  UBTC1CON127_100 U100 (O[100], I[100]);
  UBTC1CON127_101 U101 (O[101], I[101]);
  UBTC1CON127_102 U102 (O[102], I[102]);
  UBTC1CON127_103 U103 (O[103], I[103]);
  UBTC1CON127_104 U104 (O[104], I[104]);
  UBTC1CON127_105 U105 (O[105], I[105]);
  UBTC1CON127_106 U106 (O[106], I[106]);
  UBTC1CON127_107 U107 (O[107], I[107]);
  UBTC1CON127_108 U108 (O[108], I[108]);
  UBTC1CON127_109 U109 (O[109], I[109]);
  UBTC1CON127_110 U110 (O[110], I[110]);
  UBTC1CON127_111 U111 (O[111], I[111]);
  UBTC1CON127_112 U112 (O[112], I[112]);
  UBTC1CON127_113 U113 (O[113], I[113]);
  UBTC1CON127_114 U114 (O[114], I[114]);
  UBTC1CON127_115 U115 (O[115], I[115]);
  UBTC1CON127_116 U116 (O[116], I[116]);
  UBTC1CON127_117 U117 (O[117], I[117]);
  UBTC1CON127_118 U118 (O[118], I[118]);
  UBTC1CON127_119 U119 (O[119], I[119]);
  UBTC1CON127_120 U120 (O[120], I[120]);
  UBTC1CON127_121 U121 (O[121], I[121]);
  UBTC1CON127_122 U122 (O[122], I[122]);
  UBTC1CON127_123 U123 (O[123], I[123]);
  UBTC1CON127_124 U124 (O[124], I[124]);
  UBTC1CON127_125 U125 (O[125], I[125]);
  UBTC1CON127_126 U126 (O[126], I[126]);
  UBTCTCONV_127_127 U127 (O[127], I[127]);
endmodule

