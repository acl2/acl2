
module top;
wire foo;
if (0)
  begin : foo
  end
else
  begin: bar
  end

endmodule
