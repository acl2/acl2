// SV - Symbolic Vector Hardware Analysis Framework
// Copyright (C) 2014-2015 Centaur Technology
//
// Contact:
//   Centaur Technology Formal Verification Group
//   7600-C N. Capital of Texas Highway, Suite 300, Austin, TX 78731, USA.
//   http://www.centtech.com/
//
// License: (An MIT/X11-style license)
//
//   Permission is hereby granted, free of charge, to any person obtaining a
//   copy of this software and associated documentation files (the "Software"),
//   to deal in the Software without restriction, including without limitation
//   the rights to use, copy, modify, merge, publish, distribute, sublicense,
//   and/or sell copies of the Software, and to permit persons to whom the
//   Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in
//   all copies or substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//   FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//   DEALINGS IN THE SOFTWARE.
//
// Original author: Sol Swords <sswords@centtech.com>

function automatic [31:0] maj (logic [31:0] a, b, c);
  maj = (a & b) | (b & c) | (a & c);
endfunction // maj

function automatic [31:0] sum (logic [31:0] a, b, c);
  sum = a ^ b ^ c;
endfunction // sum

function automatic [31:0] sum4 (logic [31:0] a, b, c, d);
  sum4 = sum(d, sum(c, b, a), maj(c, b, a));
endfunction

function automatic [31:0] maj4 (logic [31:0] a, b, c, d);
  maj4 = maj(d, sum(c, b, a), maj(c, b, a));
endfunction



module spec (input logic [127:0] in,
	     output [127:0] out);

  logic [31:0] a, b, c, d;
   assign {a, b, c, d} = in;

   assign out = { sum4(a, b, c, d), maj4(a, b, c, d) };

endmodule // spec
 
